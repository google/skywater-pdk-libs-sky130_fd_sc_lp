* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
X0 a_202_119# a_407_93# a_56_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_978_67# a_840_95# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1273_137# a_978_67# a_1375_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND SCE a_407_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1840_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_2714_451# a_1840_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 a_1273_137# a_840_95# a_1359_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_2574_119# a_2211_428# a_2415_137# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 VPWR SCE a_245_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_323_119# a_407_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1840_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND SET_B a_2574_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_124_119# SCE a_202_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1670_93# a_1273_137# a_1423_401# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 VPWR SET_B a_2415_137# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 a_3289_47# a_2415_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_245_481# D a_202_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_978_67# a_840_95# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_2116_119# a_840_95# a_2211_428# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 VGND a_3289_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VGND SET_B a_1670_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 VPWR a_2415_137# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_2211_428# a_978_67# a_2367_163# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 Q a_3289_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_1796_379# a_1840_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 a_202_119# a_978_67# a_1273_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR SCE a_407_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_2211_428# a_840_95# a_2313_506# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VGND a_1423_401# a_2116_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X29 a_2415_137# a_2211_428# a_2714_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X30 a_3289_47# a_2415_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 VGND a_2415_137# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_1375_463# a_1423_401# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_2313_506# a_2415_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 a_2415_137# a_1840_21# a_2574_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 VPWR CLK_N a_840_95# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 a_202_119# D a_323_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_2367_163# a_2415_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 VPWR a_3289_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 Q_N a_2415_137# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X40 VPWR SET_B a_1423_401# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X41 Q_N a_2415_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X42 a_202_119# a_840_95# a_1273_137# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X43 a_1359_137# a_1423_401# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_1423_401# a_1840_21# a_1670_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X45 a_1423_401# a_1273_137# a_1796_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X46 a_56_481# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X47 VPWR a_1423_401# a_2116_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X48 Q a_3289_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X49 VGND SCD a_124_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X50 a_2116_379# a_978_67# a_2211_428# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X51 VGND CLK_N a_840_95# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
