* File: sky130_fd_sc_lp__iso0n_lp.pxi.spice
* Created: Fri Aug 28 10:40:34 2020
* 
x_PM_SKY130_FD_SC_LP__ISO0N_LP%A N_A_M1009_g N_A_M1007_g N_A_M1005_g A
+ N_A_c_49_n N_A_c_50_n PM_SKY130_FD_SC_LP__ISO0N_LP%A
x_PM_SKY130_FD_SC_LP__ISO0N_LP%SLEEP_B N_SLEEP_B_M1008_g N_SLEEP_B_M1000_g
+ N_SLEEP_B_M1001_g SLEEP_B N_SLEEP_B_c_85_n N_SLEEP_B_c_88_n
+ PM_SKY130_FD_SC_LP__ISO0N_LP%SLEEP_B
x_PM_SKY130_FD_SC_LP__ISO0N_LP%A_138_93# N_A_138_93#_M1007_s N_A_138_93#_M1005_d
+ N_A_138_93#_c_124_n N_A_138_93#_M1002_g N_A_138_93#_M1003_g
+ N_A_138_93#_c_125_n N_A_138_93#_M1004_g N_A_138_93#_M1006_g
+ N_A_138_93#_c_126_n N_A_138_93#_c_127_n N_A_138_93#_c_128_n
+ N_A_138_93#_c_144_n N_A_138_93#_c_134_n N_A_138_93#_c_135_n
+ N_A_138_93#_c_129_n N_A_138_93#_c_130_n N_A_138_93#_c_131_n
+ PM_SKY130_FD_SC_LP__ISO0N_LP%A_138_93#
x_PM_SKY130_FD_SC_LP__ISO0N_LP%VPWR N_VPWR_M1009_s N_VPWR_M1001_d N_VPWR_c_198_n
+ N_VPWR_c_199_n N_VPWR_c_200_n N_VPWR_c_201_n VPWR N_VPWR_c_202_n
+ N_VPWR_c_203_n N_VPWR_c_197_n N_VPWR_c_205_n VPWR
+ PM_SKY130_FD_SC_LP__ISO0N_LP%VPWR
x_PM_SKY130_FD_SC_LP__ISO0N_LP%X N_X_M1004_d N_X_M1006_d X X X X X N_X_c_233_n X
+ X X X X PM_SKY130_FD_SC_LP__ISO0N_LP%X
x_PM_SKY130_FD_SC_LP__ISO0N_LP%KAGND N_KAGND_M1008_d KAGND N_KAGND_c_247_n KAGND
+ PM_SKY130_FD_SC_LP__ISO0N_LP%KAGND
x_PM_SKY130_FD_SC_LP__ISO0N_LP%VGND VGND N_VGND_c_272_n N_VGND_c_273_n VGND
+ PM_SKY130_FD_SC_LP__ISO0N_LP%VGND
cc_1 VNB N_A_M1009_g 4.91509e-19 $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.655
cc_2 VNB N_A_M1007_g 0.04066f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.675
cc_3 VNB N_A_M1005_g 4.04224e-19 $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=2.655
cc_4 VNB N_A_c_49_n 0.0113041f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.48
cc_5 VNB N_A_c_50_n 0.0729266f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.48
cc_6 VNB N_SLEEP_B_M1008_g 0.0427862f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.655
cc_7 VNB N_SLEEP_B_M1000_g 3.53996e-19 $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.675
cc_8 VNB N_SLEEP_B_M1001_g 3.97322e-19 $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=2.655
cc_9 VNB N_SLEEP_B_c_85_n 0.0544878f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.48
cc_10 VNB N_A_138_93#_c_124_n 0.0216814f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.675
cc_11 VNB N_A_138_93#_c_125_n 0.0198956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_138_93#_c_126_n 0.0179657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_138_93#_c_127_n 0.0331499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_138_93#_c_128_n 0.00947454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_138_93#_c_129_n 6.61939e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_138_93#_c_130_n 0.00637441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_138_93#_c_131_n 0.0672542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_197_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_X_c_233_n 0.0627826f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.48
cc_20 VNB N_KAGND_c_247_n 0.00995849f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=0.675
cc_21 VNB KAGND 0.0518763f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.48
cc_22 VNB N_VGND_c_272_n 0.10078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_273_n 0.209029f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.645
cc_24 VPB N_A_M1009_g 0.0707471f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.655
cc_25 VPB N_A_M1005_g 0.0463725f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=2.655
cc_26 VPB N_A_c_49_n 0.0211409f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.48
cc_27 VPB N_SLEEP_B_M1000_g 0.0451068f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=0.675
cc_28 VPB N_SLEEP_B_M1001_g 0.0511816f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=2.655
cc_29 VPB N_SLEEP_B_c_88_n 0.00506395f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.48
cc_30 VPB N_A_138_93#_M1003_g 0.018301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_138_93#_M1006_g 0.0203789f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.48
cc_32 VPB N_A_138_93#_c_134_n 0.0158972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_A_138_93#_c_135_n 0.00907651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_138_93#_c_130_n 0.00185311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_138_93#_c_131_n 0.00278135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_198_n 0.0340105f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.645
cc_37 VPB N_VPWR_c_199_n 0.012785f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_38 VPB N_VPWR_c_200_n 0.0113717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_201_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.48
cc_40 VPB N_VPWR_c_202_n 0.041662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_203_n 0.0200089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_197_n 0.0865823f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_205_n 0.0101318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_X_c_233_n 0.0680606f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.48
cc_45 N_A_M1007_g N_SLEEP_B_M1008_g 0.0429872f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_46 N_A_M1005_g N_SLEEP_B_M1000_g 0.0447736f $X=1.03 $Y=2.655 $X2=0 $Y2=0
cc_47 N_A_c_49_n N_SLEEP_B_c_85_n 9.69581e-19 $X=0.87 $Y=1.48 $X2=0 $Y2=0
cc_48 N_A_c_50_n N_SLEEP_B_c_85_n 0.0429872f $X=1.03 $Y=1.48 $X2=0 $Y2=0
cc_49 N_A_M1005_g N_SLEEP_B_c_88_n 6.98642e-19 $X=1.03 $Y=2.655 $X2=0 $Y2=0
cc_50 N_A_c_49_n N_SLEEP_B_c_88_n 0.0242136f $X=0.87 $Y=1.48 $X2=0 $Y2=0
cc_51 N_A_c_50_n N_SLEEP_B_c_88_n 0.0010167f $X=1.03 $Y=1.48 $X2=0 $Y2=0
cc_52 N_A_M1007_g N_A_138_93#_c_126_n 0.0122756f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_53 N_A_M1007_g N_A_138_93#_c_127_n 0.00808815f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_54 N_A_c_49_n N_A_138_93#_c_127_n 0.00783665f $X=0.87 $Y=1.48 $X2=0 $Y2=0
cc_55 N_A_M1007_g N_A_138_93#_c_128_n 0.00418238f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_56 N_A_c_49_n N_A_138_93#_c_128_n 0.0281058f $X=0.87 $Y=1.48 $X2=0 $Y2=0
cc_57 N_A_c_50_n N_A_138_93#_c_128_n 0.00900675f $X=1.03 $Y=1.48 $X2=0 $Y2=0
cc_58 N_A_M1009_g N_A_138_93#_c_144_n 0.00272577f $X=0.67 $Y=2.655 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_A_138_93#_c_144_n 0.0158236f $X=1.03 $Y=2.655 $X2=0 $Y2=0
cc_60 N_A_M1009_g N_A_138_93#_c_135_n 8.4399e-19 $X=0.67 $Y=2.655 $X2=0 $Y2=0
cc_61 N_A_M1005_g N_A_138_93#_c_135_n 0.00615374f $X=1.03 $Y=2.655 $X2=0 $Y2=0
cc_62 N_A_c_49_n N_A_138_93#_c_135_n 6.23937e-19 $X=0.87 $Y=1.48 $X2=0 $Y2=0
cc_63 N_A_M1009_g N_VPWR_c_198_n 0.0129354f $X=0.67 $Y=2.655 $X2=0 $Y2=0
cc_64 N_A_M1005_g N_VPWR_c_198_n 0.00177594f $X=1.03 $Y=2.655 $X2=0 $Y2=0
cc_65 N_A_M1009_g N_VPWR_c_202_n 0.00424179f $X=0.67 $Y=2.655 $X2=0 $Y2=0
cc_66 N_A_M1005_g N_VPWR_c_202_n 0.00489592f $X=1.03 $Y=2.655 $X2=0 $Y2=0
cc_67 N_A_M1009_g N_VPWR_c_197_n 0.0043341f $X=0.67 $Y=2.655 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_VPWR_c_197_n 0.00515964f $X=1.03 $Y=2.655 $X2=0 $Y2=0
cc_69 N_A_M1007_g N_KAGND_c_247_n 0.00187745f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_70 N_A_M1007_g KAGND 0.00411914f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_71 N_A_M1007_g N_VGND_c_272_n 0.00489592f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_72 N_A_M1007_g N_VGND_c_273_n 0.00310524f $X=1.03 $Y=0.675 $X2=0 $Y2=0
cc_73 N_SLEEP_B_M1008_g N_A_138_93#_c_126_n 0.00205686f $X=1.39 $Y=0.675 $X2=0
+ $Y2=0
cc_74 N_SLEEP_B_M1008_g N_A_138_93#_c_127_n 0.012803f $X=1.39 $Y=0.675 $X2=0
+ $Y2=0
cc_75 N_SLEEP_B_c_85_n N_A_138_93#_c_127_n 0.0145449f $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_76 N_SLEEP_B_c_88_n N_A_138_93#_c_127_n 0.0501725f $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_77 N_SLEEP_B_M1000_g N_A_138_93#_c_144_n 0.0165672f $X=1.46 $Y=2.655 $X2=0
+ $Y2=0
cc_78 N_SLEEP_B_M1001_g N_A_138_93#_c_144_n 0.00237248f $X=1.82 $Y=2.655 $X2=0
+ $Y2=0
cc_79 N_SLEEP_B_M1000_g N_A_138_93#_c_134_n 0.0108452f $X=1.46 $Y=2.655 $X2=0
+ $Y2=0
cc_80 N_SLEEP_B_M1001_g N_A_138_93#_c_134_n 0.0154529f $X=1.82 $Y=2.655 $X2=0
+ $Y2=0
cc_81 N_SLEEP_B_c_85_n N_A_138_93#_c_134_n 6.30592e-19 $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_82 N_SLEEP_B_c_88_n N_A_138_93#_c_134_n 0.0380418f $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_83 N_SLEEP_B_M1000_g N_A_138_93#_c_135_n 0.00278249f $X=1.46 $Y=2.655 $X2=0
+ $Y2=0
cc_84 N_SLEEP_B_c_85_n N_A_138_93#_c_135_n 4.151e-19 $X=1.82 $Y=1.48 $X2=0 $Y2=0
cc_85 N_SLEEP_B_c_88_n N_A_138_93#_c_135_n 0.00712997f $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_86 N_SLEEP_B_M1001_g N_A_138_93#_c_130_n 0.00247387f $X=1.82 $Y=2.655 $X2=0
+ $Y2=0
cc_87 N_SLEEP_B_c_85_n N_A_138_93#_c_130_n 0.00379155f $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_88 N_SLEEP_B_c_88_n N_A_138_93#_c_130_n 0.0207142f $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_89 N_SLEEP_B_M1001_g N_A_138_93#_c_131_n 0.0250748f $X=1.82 $Y=2.655 $X2=0
+ $Y2=0
cc_90 N_SLEEP_B_c_85_n N_A_138_93#_c_131_n 0.0123594f $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_91 N_SLEEP_B_c_88_n N_A_138_93#_c_131_n 7.59611e-19 $X=1.82 $Y=1.48 $X2=0
+ $Y2=0
cc_92 N_SLEEP_B_M1001_g N_VPWR_c_199_n 0.0136826f $X=1.82 $Y=2.655 $X2=0 $Y2=0
cc_93 N_SLEEP_B_M1000_g N_VPWR_c_202_n 0.00489592f $X=1.46 $Y=2.655 $X2=0 $Y2=0
cc_94 N_SLEEP_B_M1001_g N_VPWR_c_202_n 0.00510437f $X=1.82 $Y=2.655 $X2=0 $Y2=0
cc_95 N_SLEEP_B_M1000_g N_VPWR_c_197_n 0.00515964f $X=1.46 $Y=2.655 $X2=0 $Y2=0
cc_96 N_SLEEP_B_M1001_g N_VPWR_c_197_n 0.00515964f $X=1.82 $Y=2.655 $X2=0 $Y2=0
cc_97 N_SLEEP_B_M1008_g N_KAGND_c_247_n 0.00981164f $X=1.39 $Y=0.675 $X2=0 $Y2=0
cc_98 N_SLEEP_B_M1008_g KAGND 0.00339751f $X=1.39 $Y=0.675 $X2=0 $Y2=0
cc_99 N_SLEEP_B_M1008_g N_VGND_c_272_n 0.00487685f $X=1.39 $Y=0.675 $X2=0 $Y2=0
cc_100 N_SLEEP_B_M1008_g N_VGND_c_273_n 0.00310524f $X=1.39 $Y=0.675 $X2=0 $Y2=0
cc_101 N_A_138_93#_c_134_n N_VPWR_M1001_d 0.0107054f $X=2.275 $Y=2.04 $X2=0
+ $Y2=0
cc_102 N_A_138_93#_c_144_n N_VPWR_c_198_n 0.0110409f $X=1.245 $Y=2.655 $X2=0
+ $Y2=0
cc_103 N_A_138_93#_M1003_g N_VPWR_c_199_n 0.0295377f $X=2.39 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_A_138_93#_M1006_g N_VPWR_c_199_n 0.00628811f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_A_138_93#_c_144_n N_VPWR_c_199_n 0.0167476f $X=1.245 $Y=2.655 $X2=0
+ $Y2=0
cc_106 N_A_138_93#_c_134_n N_VPWR_c_199_n 0.0432166f $X=2.275 $Y=2.04 $X2=0
+ $Y2=0
cc_107 N_A_138_93#_c_144_n N_VPWR_c_202_n 0.0070281f $X=1.245 $Y=2.655 $X2=0
+ $Y2=0
cc_108 N_A_138_93#_M1006_g N_VPWR_c_203_n 0.00583607f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_A_138_93#_M1006_g N_VPWR_c_197_n 0.0114293f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_138_93#_c_144_n N_VPWR_c_197_n 0.0108177f $X=1.245 $Y=2.655 $X2=0
+ $Y2=0
cc_111 N_A_138_93#_c_134_n A_493_367# 0.00106236f $X=2.275 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_138_93#_c_125_n N_X_c_233_n 0.0341466f $X=2.75 $Y=1.005 $X2=0 $Y2=0
cc_113 N_A_138_93#_c_129_n N_X_c_233_n 0.0145272f $X=2.48 $Y=1.225 $X2=0 $Y2=0
cc_114 N_A_138_93#_c_130_n N_X_c_233_n 0.0544779f $X=2.48 $Y=1.955 $X2=0 $Y2=0
cc_115 N_A_138_93#_c_124_n N_KAGND_c_247_n 0.00440396f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_116 N_A_138_93#_c_126_n N_KAGND_c_247_n 0.00891849f $X=0.815 $Y=0.675 $X2=0
+ $Y2=0
cc_117 N_A_138_93#_c_127_n N_KAGND_c_247_n 0.0490124f $X=2.275 $Y=1.14 $X2=0
+ $Y2=0
cc_118 N_A_138_93#_c_124_n KAGND 0.00500783f $X=2.39 $Y=1.17 $X2=0 $Y2=0
cc_119 N_A_138_93#_c_125_n KAGND 0.00972074f $X=2.75 $Y=1.005 $X2=0 $Y2=0
cc_120 N_A_138_93#_c_126_n KAGND 0.0342324f $X=0.815 $Y=0.675 $X2=0 $Y2=0
cc_121 N_A_138_93#_c_127_n KAGND 0.0202587f $X=2.275 $Y=1.14 $X2=0 $Y2=0
cc_122 N_A_138_93#_c_129_n KAGND 0.0161286f $X=2.48 $Y=1.225 $X2=0 $Y2=0
cc_123 N_A_138_93#_c_131_n KAGND 7.95231e-19 $X=2.515 $Y=1.17 $X2=0 $Y2=0
cc_124 N_A_138_93#_c_124_n N_VGND_c_272_n 0.00510437f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_125 N_A_138_93#_c_125_n N_VGND_c_272_n 0.00510437f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_126 N_A_138_93#_c_126_n N_VGND_c_272_n 0.00841458f $X=0.815 $Y=0.675 $X2=0
+ $Y2=0
cc_127 N_A_138_93#_c_124_n N_VGND_c_273_n 0.00310524f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_128 N_A_138_93#_c_125_n N_VGND_c_273_n 0.00310524f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_129 N_A_138_93#_c_126_n N_VGND_c_273_n 0.00145903f $X=0.815 $Y=0.675 $X2=0
+ $Y2=0
cc_130 N_VPWR_c_199_n A_493_367# 0.00103544f $X=2.175 $Y=2.38 $X2=-0.19
+ $Y2=-0.245
cc_131 N_VPWR_c_197_n N_X_M1006_d 0.00319521f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_132 N_VPWR_c_203_n N_X_c_233_n 0.0287379f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_133 N_VPWR_c_197_n N_X_c_233_n 0.0162509f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_134 N_X_c_233_n N_KAGND_c_247_n 0.0019229f $X=2.965 $Y=0.72 $X2=0 $Y2=0
cc_135 N_X_M1004_d KAGND 0.00111628f $X=2.825 $Y=0.465 $X2=0 $Y2=0
cc_136 N_X_c_233_n KAGND 0.0443903f $X=2.965 $Y=0.72 $X2=0 $Y2=0
cc_137 N_X_c_233_n N_VGND_c_272_n 0.0128756f $X=2.965 $Y=0.72 $X2=0 $Y2=0
cc_138 N_X_c_233_n N_VGND_c_273_n 0.00192863f $X=2.965 $Y=0.72 $X2=0 $Y2=0
cc_139 A_221_93# KAGND 0.00225912f $X=1.105 $Y=0.465 $X2=2.16 $Y2=0.558
cc_140 KAGND A_493_93# 0.00225631f $X=2.16 $Y=0.558 $X2=-0.19 $Y2=-0.245
cc_141 N_KAGND_c_247_n N_VGND_c_272_n 0.0310195f $X=2.11 $Y=0.555 $X2=0 $Y2=0
cc_142 KAGND N_VGND_c_272_n 0.0117374f $X=2.16 $Y=0.558 $X2=0 $Y2=0
cc_143 N_KAGND_c_247_n N_VGND_c_273_n 0.00876018f $X=2.11 $Y=0.555 $X2=0 $Y2=0
cc_144 KAGND N_VGND_c_273_n 0.298194f $X=2.16 $Y=0.558 $X2=0 $Y2=0
