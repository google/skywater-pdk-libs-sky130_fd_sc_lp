* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
X0 a_367_491# a_215_62# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_748_47# a_758_359# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_758_359# a_1266_147# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VGND a_1266_147# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_608_491# a_367_491# a_713_491# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR GATE a_215_62# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_608_491# a_215_62# a_748_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_713_491# a_758_359# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_536_491# a_215_62# a_608_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_46_62# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_46_62# a_568_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 Q a_758_359# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_46_62# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 Q a_758_359# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR a_1266_147# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND GATE a_215_62# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_608_491# a_758_359# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR a_46_62# a_536_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_367_491# a_215_62# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_568_47# a_367_491# a_608_491# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_608_491# a_758_359# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND a_758_359# a_1266_147# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
