# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 1.170000 1.315000 1.390000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.295000 1.815000 7.535000 1.985000 ;
        RECT 6.295000 1.985000 6.525000 3.075000 ;
        RECT 6.485000 0.255000 6.675000 1.075000 ;
        RECT 6.485000 1.075000 7.535000 1.245000 ;
        RECT 7.195000 1.985000 7.535000 3.075000 ;
        RECT 7.345000 0.255000 7.535000 1.075000 ;
        RECT 7.355000 1.245000 7.535000 1.815000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.400000 1.365000 3.850000 1.760000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.550000  0.085000 0.890000 0.660000 ;
        RECT 2.685000  0.085000 2.945000 0.780000 ;
        RECT 4.675000  0.085000 5.005000 0.455000 ;
        RECT 5.985000  0.085000 6.315000 0.895000 ;
        RECT 6.845000  0.085000 7.175000 0.905000 ;
        RECT 7.740000  0.085000 8.035000 1.095000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.605000 2.970000 0.935000 3.245000 ;
        RECT 2.525000 2.620000 2.855000 3.245000 ;
        RECT 4.840000 2.850000 5.170000 3.245000 ;
        RECT 5.795000 2.850000 6.125000 3.245000 ;
        RECT 6.695000 2.165000 7.025000 3.245000 ;
        RECT 7.705000 1.815000 7.955000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.255000 0.380000 0.830000 ;
      RECT 0.095000 0.830000 1.230000 1.000000 ;
      RECT 0.095000 1.000000 0.450000 1.095000 ;
      RECT 0.095000 1.095000 0.265000 1.900000 ;
      RECT 0.095000 1.900000 0.425000 2.630000 ;
      RECT 0.095000 2.630000 1.285000 2.800000 ;
      RECT 0.095000 2.800000 0.435000 3.075000 ;
      RECT 0.435000 1.345000 0.685000 1.560000 ;
      RECT 0.435000 1.560000 1.655000 1.730000 ;
      RECT 1.035000 1.730000 1.205000 2.280000 ;
      RECT 1.035000 2.280000 1.840000 2.450000 ;
      RECT 1.060000 0.265000 2.515000 0.435000 ;
      RECT 1.060000 0.435000 1.230000 0.830000 ;
      RECT 1.115000 2.800000 1.285000 2.905000 ;
      RECT 1.115000 2.905000 2.190000 3.075000 ;
      RECT 1.385000 1.900000 2.165000 1.930000 ;
      RECT 1.385000 1.930000 3.695000 2.110000 ;
      RECT 1.485000 0.605000 1.930000 0.845000 ;
      RECT 1.485000 0.845000 1.655000 1.560000 ;
      RECT 1.510000 2.450000 1.840000 2.735000 ;
      RECT 1.835000 1.015000 2.165000 1.900000 ;
      RECT 2.020000 2.280000 3.195000 2.450000 ;
      RECT 2.020000 2.450000 2.190000 2.905000 ;
      RECT 2.345000 0.435000 2.515000 1.015000 ;
      RECT 2.345000 1.015000 2.705000 1.265000 ;
      RECT 2.345000 1.475000 3.230000 1.760000 ;
      RECT 2.920000 0.965000 4.530000 1.195000 ;
      RECT 2.920000 1.195000 3.230000 1.475000 ;
      RECT 3.025000 2.450000 3.195000 2.765000 ;
      RECT 3.025000 2.765000 4.540000 3.075000 ;
      RECT 3.115000 0.465000 3.375000 0.625000 ;
      RECT 3.115000 0.625000 5.080000 0.795000 ;
      RECT 3.365000 2.110000 3.695000 2.160000 ;
      RECT 3.365000 2.160000 5.080000 2.340000 ;
      RECT 3.365000 2.340000 3.635000 2.535000 ;
      RECT 3.805000 2.510000 5.975000 2.680000 ;
      RECT 3.805000 2.680000 4.540000 2.765000 ;
      RECT 4.200000 1.195000 4.530000 1.990000 ;
      RECT 4.700000 0.795000 5.080000 2.160000 ;
      RECT 5.250000 1.065000 6.315000 1.235000 ;
      RECT 5.250000 1.235000 5.420000 2.010000 ;
      RECT 5.250000 2.010000 5.625000 2.340000 ;
      RECT 5.465000 0.255000 5.795000 1.065000 ;
      RECT 5.600000 1.405000 5.975000 1.665000 ;
      RECT 5.795000 1.665000 5.975000 2.510000 ;
      RECT 6.145000 1.235000 6.315000 1.415000 ;
      RECT 6.145000 1.415000 7.155000 1.585000 ;
  END
END sky130_fd_sc_lp__dlclkp_4
