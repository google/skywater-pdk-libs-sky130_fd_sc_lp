# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21boi_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a21boi_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.460000 1.315000 1.790000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.810000 0.835000 1.140000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.825000 2.855000 1.495000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 0.265000 1.665000 0.675000 ;
        RECT 1.495000 0.675000 1.665000 1.920000 ;
        RECT 1.495000 1.920000 1.865000 2.025000 ;
        RECT 1.495000 2.025000 2.045000 2.150000 ;
        RECT 1.695000 2.150000 2.045000 3.065000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.125000  2.025000 0.455000 2.330000 ;
      RECT 0.125000  2.330000 1.515000 2.500000 ;
      RECT 0.125000  2.500000 0.455000 3.065000 ;
      RECT 0.405000  0.085000 0.735000 0.630000 ;
      RECT 0.655000  2.680000 0.985000 3.245000 ;
      RECT 1.185000  2.500000 1.515000 3.065000 ;
      RECT 1.845000  1.070000 2.215000 1.675000 ;
      RECT 1.845000  1.675000 3.230000 1.740000 ;
      RECT 2.015000  0.085000 2.345000 0.675000 ;
      RECT 2.045000  1.740000 3.230000 1.845000 ;
      RECT 2.370000  2.025000 2.700000 3.245000 ;
      RECT 2.900000  0.265000 3.230000 0.645000 ;
      RECT 2.900000  1.845000 3.230000 3.065000 ;
      RECT 3.060000  0.645000 3.230000 1.675000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__a21boi_lp
END LIBRARY
