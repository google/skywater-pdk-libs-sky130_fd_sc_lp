* NGSPICE file created from sky130_fd_sc_lp__and2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and2b_1 A_N B VGND VNB VPB VPWR X
M1000 a_217_131# a_27_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.701e+11p pd=1.65e+06u as=5.817e+11p ps=5.07e+06u
M1001 VPWR B a_217_131# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_217_131# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1003 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=4.053e+11p pd=3.92e+06u as=1.113e+11p ps=1.37e+06u
M1004 VGND B a_300_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 X a_217_131# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1006 a_300_131# a_27_47# a_217_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VPWR A_N a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

