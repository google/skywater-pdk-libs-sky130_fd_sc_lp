* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__clkinvlp_16 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VGND A a_426_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X3 VGND A a_1058_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 Y A a_1216_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_900_67# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_268_67# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_584_67# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X13 VGND A a_742_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X14 a_1058_67# A Y VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_742_67# A Y VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X17 a_1374_67# A Y VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 Y A a_900_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X21 Y A a_1532_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X22 a_110_67# A Y VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X23 a_1532_67# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 VGND A a_110_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X26 a_426_67# A Y VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X29 Y A a_584_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X30 a_1216_67# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X31 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 VGND A a_1374_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X34 Y A a_268_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
