* NGSPICE file created from sky130_fd_sc_lp__nor4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
M1000 Y a_80_131# a_451_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.78e+11p pd=3.12e+06u as=4.914e+11p ps=3.3e+06u
M1001 a_271_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=3.864e+11p ps=3.3e+06u
M1002 VGND B Y VNB nshort w=840000u l=150000u
+  ad=8.211e+11p pd=7.12e+06u as=5.082e+11p ps=4.57e+06u
M1003 a_343_367# B a_271_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.914e+11p pd=3.3e+06u as=0p ps=0u
M1004 VGND a_80_131# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND D_N a_80_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_451_367# C a_343_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y C VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR D_N a_80_131# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

