* File: sky130_fd_sc_lp__ebufn_2.pxi.spice
* Created: Fri Aug 28 10:31:41 2020
* 
x_PM_SKY130_FD_SC_LP__EBUFN_2%A_96_21# N_A_96_21#_M1005_d N_A_96_21#_M1011_d
+ N_A_96_21#_M1001_g N_A_96_21#_M1002_g N_A_96_21#_M1010_g N_A_96_21#_M1009_g
+ N_A_96_21#_c_92_n N_A_96_21#_c_98_n N_A_96_21#_c_99_n N_A_96_21#_c_100_n
+ N_A_96_21#_c_101_n N_A_96_21#_c_102_n N_A_96_21#_c_93_n N_A_96_21#_c_104_n
+ N_A_96_21#_c_105_n N_A_96_21#_c_94_n N_A_96_21#_c_95_n
+ PM_SKY130_FD_SC_LP__EBUFN_2%A_96_21#
x_PM_SKY130_FD_SC_LP__EBUFN_2%A_284_21# N_A_284_21#_M1008_s N_A_284_21#_M1006_s
+ N_A_284_21#_c_200_n N_A_284_21#_M1004_g N_A_284_21#_c_201_n
+ N_A_284_21#_c_202_n N_A_284_21#_c_203_n N_A_284_21#_M1007_g
+ N_A_284_21#_c_204_n N_A_284_21#_c_205_n N_A_284_21#_c_206_n
+ N_A_284_21#_c_228_p N_A_284_21#_c_207_n N_A_284_21#_c_208_n
+ N_A_284_21#_c_209_n N_A_284_21#_c_210_n PM_SKY130_FD_SC_LP__EBUFN_2%A_284_21#
x_PM_SKY130_FD_SC_LP__EBUFN_2%TE_B N_TE_B_c_274_n N_TE_B_M1000_g N_TE_B_c_267_n
+ N_TE_B_c_268_n N_TE_B_c_277_n N_TE_B_M1003_g N_TE_B_c_269_n N_TE_B_M1006_g
+ N_TE_B_M1008_g N_TE_B_c_271_n TE_B TE_B N_TE_B_c_272_n N_TE_B_c_273_n
+ PM_SKY130_FD_SC_LP__EBUFN_2%TE_B
x_PM_SKY130_FD_SC_LP__EBUFN_2%A N_A_M1011_g N_A_M1005_g N_A_c_350_n N_A_c_355_n
+ A A N_A_c_351_n N_A_c_352_n PM_SKY130_FD_SC_LP__EBUFN_2%A
x_PM_SKY130_FD_SC_LP__EBUFN_2%A_39_367# N_A_39_367#_M1002_s N_A_39_367#_M1010_s
+ N_A_39_367#_M1003_d N_A_39_367#_c_385_n N_A_39_367#_c_386_n
+ N_A_39_367#_c_393_n N_A_39_367#_c_387_n N_A_39_367#_c_398_n
+ N_A_39_367#_c_388_n N_A_39_367#_c_389_n N_A_39_367#_c_403_n
+ PM_SKY130_FD_SC_LP__EBUFN_2%A_39_367#
x_PM_SKY130_FD_SC_LP__EBUFN_2%Z N_Z_M1001_d N_Z_M1002_d N_Z_c_437_n N_Z_c_438_n
+ N_Z_c_440_n N_Z_c_441_n N_Z_c_451_n N_Z_c_461_n Z Z
+ PM_SKY130_FD_SC_LP__EBUFN_2%Z
x_PM_SKY130_FD_SC_LP__EBUFN_2%VPWR N_VPWR_M1000_s N_VPWR_M1006_d N_VPWR_c_473_n
+ N_VPWR_c_474_n N_VPWR_c_475_n N_VPWR_c_476_n VPWR N_VPWR_c_477_n
+ N_VPWR_c_478_n N_VPWR_c_472_n N_VPWR_c_480_n PM_SKY130_FD_SC_LP__EBUFN_2%VPWR
x_PM_SKY130_FD_SC_LP__EBUFN_2%A_27_47# N_A_27_47#_M1001_s N_A_27_47#_M1009_s
+ N_A_27_47#_M1007_d N_A_27_47#_c_526_n N_A_27_47#_c_531_n N_A_27_47#_c_527_n
+ N_A_27_47#_c_536_n N_A_27_47#_c_537_n N_A_27_47#_c_528_n N_A_27_47#_c_529_n
+ N_A_27_47#_c_530_n PM_SKY130_FD_SC_LP__EBUFN_2%A_27_47#
x_PM_SKY130_FD_SC_LP__EBUFN_2%VGND N_VGND_M1004_s N_VGND_M1008_d N_VGND_c_575_n
+ N_VGND_c_576_n VGND N_VGND_c_577_n N_VGND_c_578_n N_VGND_c_579_n
+ N_VGND_c_580_n N_VGND_c_581_n N_VGND_c_582_n PM_SKY130_FD_SC_LP__EBUFN_2%VGND
cc_1 VNB N_A_96_21#_M1001_g 0.0255833f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.655
cc_2 VNB N_A_96_21#_M1002_g 0.00160006f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_3 VNB N_A_96_21#_M1010_g 0.00152339f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_4 VNB N_A_96_21#_M1009_g 0.0230116f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.655
cc_5 VNB N_A_96_21#_c_92_n 0.0088736f $X=-0.19 $Y=-0.245 $X2=2.315 $Y2=1.46
cc_6 VNB N_A_96_21#_c_93_n 0.024461f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=2.435
cc_7 VNB N_A_96_21#_c_94_n 0.029726f $X=-0.19 $Y=-0.245 $X2=4.035 $Y2=0.905
cc_8 VNB N_A_96_21#_c_95_n 0.0423951f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.46
cc_9 VNB N_A_284_21#_c_200_n 0.0171726f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.295
cc_10 VNB N_A_284_21#_c_201_n 0.0131969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_284_21#_c_202_n 0.00726992f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.625
cc_12 VNB N_A_284_21#_c_203_n 0.0199408f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_13 VNB N_A_284_21#_c_204_n 0.0336091f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.625
cc_14 VNB N_A_284_21#_c_205_n 0.0356991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_284_21#_c_206_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.295
cc_16 VNB N_A_284_21#_c_207_n 0.00570941f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.46
cc_17 VNB N_A_284_21#_c_208_n 0.00762634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_284_21#_c_209_n 0.0436387f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=1.625
cc_19 VNB N_A_284_21#_c_210_n 0.00356436f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=2.53
cc_20 VNB N_TE_B_c_267_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_TE_B_c_268_n 0.00559972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_TE_B_c_269_n 0.0267714f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.655
cc_23 VNB N_TE_B_M1008_g 0.0239914f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_24 VNB N_TE_B_c_271_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.295
cc_25 VNB N_TE_B_c_272_n 0.0299636f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.46
cc_26 VNB N_TE_B_c_273_n 0.00167757f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.46
cc_27 VNB N_A_M1005_g 0.0288087f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.295
cc_28 VNB N_A_c_350_n 0.013025f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.625
cc_29 VNB N_A_c_351_n 0.0168177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_c_352_n 0.00586238f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.295
cc_31 VNB N_Z_c_437_n 0.00482248f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.295
cc_32 VNB N_Z_c_438_n 0.00738541f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.655
cc_33 VNB Z 0.0273998f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.655
cc_34 VNB N_VPWR_c_472_n 0.183584f $X=-0.19 $Y=-0.245 $X2=4.035 $Y2=2.615
cc_35 VNB N_A_27_47#_c_526_n 0.0140806f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_36 VNB N_A_27_47#_c_527_n 0.00718715f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.625
cc_37 VNB N_A_27_47#_c_528_n 0.00570274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_529_n 0.00314727f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.295
cc_39 VNB N_A_27_47#_c_530_n 0.00563257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_575_n 0.00512425f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.655
cc_41 VNB N_VGND_c_576_n 0.0349587f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_42 VNB N_VGND_c_577_n 0.0409482f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_43 VNB N_VGND_c_578_n 0.0384923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_579_n 0.0203806f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=2.53
cc_45 VNB N_VGND_c_580_n 0.255736f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=2.53
cc_46 VNB N_VGND_c_581_n 0.00480536f $X=-0.19 $Y=-0.245 $X2=4 $Y2=2.755
cc_47 VNB N_VGND_c_582_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=2.53
cc_48 VPB N_A_96_21#_M1002_g 0.0232657f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_49 VPB N_A_96_21#_M1010_g 0.0200267f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_50 VPB N_A_96_21#_c_98_n 0.0176559f $X=-0.19 $Y=1.655 $X2=2.4 $Y2=2.615
cc_51 VPB N_A_96_21#_c_99_n 0.0102947f $X=-0.19 $Y=1.655 $X2=2.995 $Y2=2.7
cc_52 VPB N_A_96_21#_c_100_n 0.00422484f $X=-0.19 $Y=1.655 $X2=2.485 $Y2=2.7
cc_53 VPB N_A_96_21#_c_101_n 0.00576138f $X=-0.19 $Y=1.655 $X2=3.835 $Y2=2.53
cc_54 VPB N_A_96_21#_c_102_n 0.0196727f $X=-0.19 $Y=1.655 $X2=4.035 $Y2=2.615
cc_55 VPB N_A_96_21#_c_93_n 0.0370709f $X=-0.19 $Y=1.655 $X2=4.15 $Y2=2.435
cc_56 VPB N_A_96_21#_c_104_n 3.20284e-19 $X=-0.19 $Y=1.655 $X2=3.08 $Y2=2.53
cc_57 VPB N_A_96_21#_c_105_n 0.0151865f $X=-0.19 $Y=1.655 $X2=4.035 $Y2=2.525
cc_58 VPB N_A_284_21#_c_207_n 0.00759081f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.46
cc_59 VPB N_TE_B_c_274_n 0.0162047f $X=-0.19 $Y=1.655 $X2=3.895 $Y2=0.695
cc_60 VPB N_TE_B_c_267_n 0.00421372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_TE_B_c_268_n 0.00251798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_TE_B_c_277_n 0.0197118f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_TE_B_c_269_n 0.0404582f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.655
cc_64 VPB N_TE_B_M1006_g 0.0253024f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_65 VPB N_TE_B_c_271_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.295
cc_66 VPB N_TE_B_c_272_n 0.0280541f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.46
cc_67 VPB N_TE_B_c_273_n 0.00111101f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.46
cc_68 VPB N_A_M1011_g 0.0491006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_c_350_n 0.0109014f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.625
cc_70 VPB N_A_c_355_n 0.0167892f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_71 VPB N_A_c_352_n 0.00758542f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.295
cc_72 VPB N_A_39_367#_c_385_n 0.00719502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_39_367#_c_386_n 0.029378f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_74 VPB N_A_39_367#_c_387_n 0.00269919f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_75 VPB N_A_39_367#_c_388_n 0.00192554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_39_367#_c_389_n 0.00172323f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.655
cc_77 VPB N_Z_c_440_n 0.00461635f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.655
cc_78 VPB N_Z_c_441_n 0.00973359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB Z 0.00719786f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.655
cc_80 VPB N_VPWR_c_473_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.655
cc_81 VPB N_VPWR_c_474_n 0.0140867f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_82 VPB N_VPWR_c_475_n 0.0438543f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_83 VPB N_VPWR_c_476_n 0.00631567f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_84 VPB N_VPWR_c_477_n 0.0397154f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.655
cc_85 VPB N_VPWR_c_478_n 0.018465f $X=-0.19 $Y=1.655 $X2=3.165 $Y2=2.53
cc_86 VPB N_VPWR_c_472_n 0.0637668f $X=-0.19 $Y=1.655 $X2=4.035 $Y2=2.615
cc_87 VPB N_VPWR_c_480_n 0.00324402f $X=-0.19 $Y=1.655 $X2=4.15 $Y2=1.135
cc_88 N_A_96_21#_c_99_n N_A_284_21#_M1006_s 0.010408f $X=2.995 $Y=2.7 $X2=0
+ $Y2=0
cc_89 N_A_96_21#_M1009_g N_A_284_21#_c_200_n 0.0144781f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_90 N_A_96_21#_c_92_n N_A_284_21#_c_201_n 0.00874973f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_91 N_A_96_21#_c_92_n N_A_284_21#_c_202_n 0.00478473f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_92 N_A_96_21#_c_95_n N_A_284_21#_c_202_n 0.0144781f $X=0.995 $Y=1.46 $X2=0
+ $Y2=0
cc_93 N_A_96_21#_c_92_n N_A_284_21#_c_204_n 0.014197f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_94 N_A_96_21#_c_92_n N_A_284_21#_c_206_n 0.004228f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_95 N_A_96_21#_c_92_n N_A_284_21#_c_207_n 0.0271261f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_96 N_A_96_21#_c_98_n N_A_284_21#_c_207_n 0.060547f $X=2.4 $Y=2.615 $X2=0
+ $Y2=0
cc_97 N_A_96_21#_c_99_n N_A_284_21#_c_207_n 0.0136682f $X=2.995 $Y=2.7 $X2=0
+ $Y2=0
cc_98 N_A_96_21#_c_92_n N_TE_B_c_267_n 0.00764923f $X=2.315 $Y=1.46 $X2=0 $Y2=0
cc_99 N_A_96_21#_M1010_g N_TE_B_c_268_n 0.0243873f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_96_21#_c_92_n N_TE_B_c_268_n 0.00581178f $X=2.315 $Y=1.46 $X2=0 $Y2=0
cc_101 N_A_96_21#_c_95_n N_TE_B_c_268_n 0.00241004f $X=0.995 $Y=1.46 $X2=0 $Y2=0
cc_102 N_A_96_21#_c_98_n N_TE_B_c_277_n 0.00382744f $X=2.4 $Y=2.615 $X2=0 $Y2=0
cc_103 N_A_96_21#_c_100_n N_TE_B_c_277_n 5.46443e-19 $X=2.485 $Y=2.7 $X2=0 $Y2=0
cc_104 N_A_96_21#_c_92_n N_TE_B_c_269_n 0.0184428f $X=2.315 $Y=1.46 $X2=0 $Y2=0
cc_105 N_A_96_21#_c_98_n N_TE_B_c_269_n 0.0113471f $X=2.4 $Y=2.615 $X2=0 $Y2=0
cc_106 N_A_96_21#_c_98_n N_TE_B_M1006_g 0.00339138f $X=2.4 $Y=2.615 $X2=0 $Y2=0
cc_107 N_A_96_21#_c_99_n N_TE_B_M1006_g 0.00342807f $X=2.995 $Y=2.7 $X2=0 $Y2=0
cc_108 N_A_96_21#_c_104_n N_TE_B_M1006_g 0.0159544f $X=3.08 $Y=2.53 $X2=0 $Y2=0
cc_109 N_A_96_21#_c_92_n N_TE_B_c_271_n 0.00449494f $X=2.315 $Y=1.46 $X2=0 $Y2=0
cc_110 N_A_96_21#_c_101_n N_TE_B_c_272_n 6.29048e-19 $X=3.835 $Y=2.53 $X2=0
+ $Y2=0
cc_111 N_A_96_21#_c_101_n N_TE_B_c_273_n 0.00660564f $X=3.835 $Y=2.53 $X2=0
+ $Y2=0
cc_112 N_A_96_21#_c_104_n N_TE_B_c_273_n 0.00768035f $X=3.08 $Y=2.53 $X2=0 $Y2=0
cc_113 N_A_96_21#_c_101_n N_A_M1011_g 0.0104163f $X=3.835 $Y=2.53 $X2=0 $Y2=0
cc_114 N_A_96_21#_c_102_n N_A_M1011_g 0.00948065f $X=4.035 $Y=2.615 $X2=0 $Y2=0
cc_115 N_A_96_21#_c_93_n N_A_M1011_g 0.00887849f $X=4.15 $Y=2.435 $X2=0 $Y2=0
cc_116 N_A_96_21#_c_104_n N_A_M1011_g 5.76141e-19 $X=3.08 $Y=2.53 $X2=0 $Y2=0
cc_117 N_A_96_21#_c_105_n N_A_M1011_g 0.00373339f $X=4.035 $Y=2.525 $X2=0 $Y2=0
cc_118 N_A_96_21#_c_93_n N_A_M1005_g 0.0190728f $X=4.15 $Y=2.435 $X2=0 $Y2=0
cc_119 N_A_96_21#_c_94_n N_A_M1005_g 0.00694532f $X=4.035 $Y=0.905 $X2=0 $Y2=0
cc_120 N_A_96_21#_c_101_n N_A_c_355_n 6.44547e-19 $X=3.835 $Y=2.53 $X2=0 $Y2=0
cc_121 N_A_96_21#_c_101_n N_A_c_352_n 0.0178279f $X=3.835 $Y=2.53 $X2=0 $Y2=0
cc_122 N_A_96_21#_c_93_n N_A_c_352_n 0.064988f $X=4.15 $Y=2.435 $X2=0 $Y2=0
cc_123 N_A_96_21#_c_105_n N_A_c_352_n 0.00359627f $X=4.035 $Y=2.525 $X2=0 $Y2=0
cc_124 N_A_96_21#_c_94_n N_A_c_352_n 0.00189076f $X=4.035 $Y=0.905 $X2=0 $Y2=0
cc_125 N_A_96_21#_M1002_g N_A_39_367#_c_385_n 5.89773e-19 $X=0.555 $Y=2.465
+ $X2=0 $Y2=0
cc_126 N_A_96_21#_M1002_g N_A_39_367#_c_386_n 0.00948285f $X=0.555 $Y=2.465
+ $X2=0 $Y2=0
cc_127 N_A_96_21#_M1010_g N_A_39_367#_c_386_n 6.13901e-19 $X=0.985 $Y=2.465
+ $X2=0 $Y2=0
cc_128 N_A_96_21#_M1002_g N_A_39_367#_c_393_n 0.0105205f $X=0.555 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_96_21#_M1010_g N_A_39_367#_c_393_n 0.0105205f $X=0.985 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_96_21#_M1010_g N_A_39_367#_c_387_n 0.00236068f $X=0.985 $Y=2.465
+ $X2=0 $Y2=0
cc_131 N_A_96_21#_c_92_n N_A_39_367#_c_387_n 0.0265018f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_132 N_A_96_21#_c_95_n N_A_39_367#_c_387_n 2.69228e-19 $X=0.995 $Y=1.46 $X2=0
+ $Y2=0
cc_133 N_A_96_21#_M1002_g N_A_39_367#_c_398_n 6.58365e-19 $X=0.555 $Y=2.465
+ $X2=0 $Y2=0
cc_134 N_A_96_21#_M1010_g N_A_39_367#_c_398_n 0.0130432f $X=0.985 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_96_21#_c_92_n N_A_39_367#_c_388_n 0.035557f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_136 N_A_96_21#_c_92_n N_A_39_367#_c_389_n 0.0192431f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_137 N_A_96_21#_c_98_n N_A_39_367#_c_389_n 0.0140923f $X=2.4 $Y=2.615 $X2=0
+ $Y2=0
cc_138 N_A_96_21#_c_98_n N_A_39_367#_c_403_n 0.0478824f $X=2.4 $Y=2.615 $X2=0
+ $Y2=0
cc_139 N_A_96_21#_c_100_n N_A_39_367#_c_403_n 0.0145003f $X=2.485 $Y=2.7 $X2=0
+ $Y2=0
cc_140 N_A_96_21#_M1001_g N_Z_c_437_n 0.0150407f $X=0.555 $Y=0.655 $X2=0 $Y2=0
cc_141 N_A_96_21#_M1009_g N_Z_c_437_n 0.00363496f $X=0.995 $Y=0.655 $X2=0 $Y2=0
cc_142 N_A_96_21#_c_92_n N_Z_c_437_n 0.016831f $X=2.315 $Y=1.46 $X2=0 $Y2=0
cc_143 N_A_96_21#_c_95_n N_Z_c_437_n 0.00270745f $X=0.995 $Y=1.46 $X2=0 $Y2=0
cc_144 N_A_96_21#_M1002_g N_Z_c_440_n 0.0163408f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_96_21#_M1010_g N_Z_c_440_n 7.94117e-19 $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_96_21#_c_92_n N_Z_c_440_n 0.00969903f $X=2.315 $Y=1.46 $X2=0 $Y2=0
cc_147 N_A_96_21#_c_95_n N_Z_c_440_n 0.00246695f $X=0.995 $Y=1.46 $X2=0 $Y2=0
cc_148 N_A_96_21#_M1001_g N_Z_c_451_n 0.00946396f $X=0.555 $Y=0.655 $X2=0 $Y2=0
cc_149 N_A_96_21#_M1009_g N_Z_c_451_n 0.00419329f $X=0.995 $Y=0.655 $X2=0 $Y2=0
cc_150 N_A_96_21#_M1001_g Z 0.0223777f $X=0.555 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A_96_21#_c_92_n Z 0.0144709f $X=2.315 $Y=1.46 $X2=0 $Y2=0
cc_152 N_A_96_21#_c_101_n N_VPWR_M1006_d 0.0117955f $X=3.835 $Y=2.53 $X2=0 $Y2=0
cc_153 N_A_96_21#_c_101_n N_VPWR_c_474_n 0.0247657f $X=3.835 $Y=2.53 $X2=0 $Y2=0
cc_154 N_A_96_21#_c_99_n N_VPWR_c_475_n 0.0113897f $X=2.995 $Y=2.7 $X2=0 $Y2=0
cc_155 N_A_96_21#_c_100_n N_VPWR_c_475_n 0.00420318f $X=2.485 $Y=2.7 $X2=0 $Y2=0
cc_156 N_A_96_21#_c_101_n N_VPWR_c_475_n 0.00224723f $X=3.835 $Y=2.53 $X2=0
+ $Y2=0
cc_157 N_A_96_21#_c_104_n N_VPWR_c_475_n 0.0036221f $X=3.08 $Y=2.53 $X2=0 $Y2=0
cc_158 N_A_96_21#_M1002_g N_VPWR_c_477_n 0.00357842f $X=0.555 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_96_21#_M1010_g N_VPWR_c_477_n 0.00357842f $X=0.985 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_96_21#_c_101_n N_VPWR_c_478_n 0.00205091f $X=3.835 $Y=2.53 $X2=0
+ $Y2=0
cc_161 N_A_96_21#_c_102_n N_VPWR_c_478_n 0.0260166f $X=4.035 $Y=2.615 $X2=0
+ $Y2=0
cc_162 N_A_96_21#_M1011_d N_VPWR_c_472_n 0.00232718f $X=3.86 $Y=2.455 $X2=0
+ $Y2=0
cc_163 N_A_96_21#_M1002_g N_VPWR_c_472_n 0.00635114f $X=0.555 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_96_21#_M1010_g N_VPWR_c_472_n 0.00537652f $X=0.985 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_96_21#_c_99_n N_VPWR_c_472_n 0.0156153f $X=2.995 $Y=2.7 $X2=0 $Y2=0
cc_166 N_A_96_21#_c_100_n N_VPWR_c_472_n 0.00550847f $X=2.485 $Y=2.7 $X2=0 $Y2=0
cc_167 N_A_96_21#_c_101_n N_VPWR_c_472_n 0.00981335f $X=3.835 $Y=2.53 $X2=0
+ $Y2=0
cc_168 N_A_96_21#_c_102_n N_VPWR_c_472_n 0.0153493f $X=4.035 $Y=2.615 $X2=0
+ $Y2=0
cc_169 N_A_96_21#_c_104_n N_VPWR_c_472_n 0.00512927f $X=3.08 $Y=2.53 $X2=0 $Y2=0
cc_170 N_A_96_21#_M1001_g N_A_27_47#_c_531_n 0.0129105f $X=0.555 $Y=0.655 $X2=0
+ $Y2=0
cc_171 N_A_96_21#_M1009_g N_A_27_47#_c_531_n 0.0139717f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_172 N_A_96_21#_c_92_n N_A_27_47#_c_528_n 0.0719464f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_173 N_A_96_21#_M1009_g N_A_27_47#_c_529_n 0.00108019f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_174 N_A_96_21#_c_92_n N_A_27_47#_c_529_n 0.0289763f $X=2.315 $Y=1.46 $X2=0
+ $Y2=0
cc_175 N_A_96_21#_c_94_n N_VGND_c_576_n 0.0191097f $X=4.035 $Y=0.905 $X2=0 $Y2=0
cc_176 N_A_96_21#_M1001_g N_VGND_c_577_n 0.00357877f $X=0.555 $Y=0.655 $X2=0
+ $Y2=0
cc_177 N_A_96_21#_M1009_g N_VGND_c_577_n 0.00357877f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_178 N_A_96_21#_c_94_n N_VGND_c_579_n 0.00662032f $X=4.035 $Y=0.905 $X2=0
+ $Y2=0
cc_179 N_A_96_21#_M1001_g N_VGND_c_580_n 0.00652668f $X=0.555 $Y=0.655 $X2=0
+ $Y2=0
cc_180 N_A_96_21#_M1009_g N_VGND_c_580_n 0.00564902f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_181 N_A_96_21#_c_94_n N_VGND_c_580_n 0.0105622f $X=4.035 $Y=0.905 $X2=0 $Y2=0
cc_182 N_A_284_21#_c_201_n N_TE_B_c_267_n 0.0187271f $X=1.92 $Y=1.26 $X2=0 $Y2=0
cc_183 N_A_284_21#_c_202_n N_TE_B_c_268_n 0.0187271f $X=1.57 $Y=1.26 $X2=0 $Y2=0
cc_184 N_A_284_21#_c_204_n N_TE_B_c_269_n 0.0187271f $X=2.605 $Y=1.26 $X2=0
+ $Y2=0
cc_185 N_A_284_21#_c_207_n N_TE_B_c_269_n 0.0131944f $X=2.74 $Y=2.28 $X2=0 $Y2=0
cc_186 N_A_284_21#_c_210_n N_TE_B_c_269_n 0.00573077f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_187 N_A_284_21#_c_205_n N_TE_B_M1008_g 0.0134967f $X=2.68 $Y=1.185 $X2=0
+ $Y2=0
cc_188 N_A_284_21#_c_228_p N_TE_B_M1008_g 0.00545376f $X=2.927 $Y=0.863 $X2=0
+ $Y2=0
cc_189 N_A_284_21#_c_207_n N_TE_B_M1008_g 0.0029973f $X=2.74 $Y=2.28 $X2=0 $Y2=0
cc_190 N_A_284_21#_c_208_n N_TE_B_M1008_g 8.98453e-19 $X=2.77 $Y=0.42 $X2=0
+ $Y2=0
cc_191 N_A_284_21#_c_209_n N_TE_B_M1008_g 0.00109563f $X=2.77 $Y=0.42 $X2=0
+ $Y2=0
cc_192 N_A_284_21#_c_210_n N_TE_B_M1008_g 0.00345432f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_193 N_A_284_21#_c_206_n N_TE_B_c_271_n 0.0187271f $X=1.995 $Y=1.26 $X2=0
+ $Y2=0
cc_194 N_A_284_21#_c_204_n N_TE_B_c_272_n 0.00158731f $X=2.605 $Y=1.26 $X2=0
+ $Y2=0
cc_195 N_A_284_21#_c_207_n N_TE_B_c_272_n 0.0245801f $X=2.74 $Y=2.28 $X2=0 $Y2=0
cc_196 N_A_284_21#_c_210_n N_TE_B_c_272_n 0.00140009f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_197 N_A_284_21#_c_207_n N_TE_B_c_273_n 0.0628885f $X=2.74 $Y=2.28 $X2=0 $Y2=0
cc_198 N_A_284_21#_c_210_n N_TE_B_c_273_n 0.0179903f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_199 N_A_284_21#_c_202_n N_A_39_367#_c_388_n 3.75348e-19 $X=1.57 $Y=1.26 $X2=0
+ $Y2=0
cc_200 N_A_284_21#_c_206_n N_A_39_367#_c_389_n 2.41418e-19 $X=1.995 $Y=1.26
+ $X2=0 $Y2=0
cc_201 N_A_284_21#_c_200_n N_A_27_47#_c_536_n 0.00199024f $X=1.495 $Y=1.185
+ $X2=0 $Y2=0
cc_202 N_A_284_21#_c_200_n N_A_27_47#_c_537_n 0.00840415f $X=1.495 $Y=1.185
+ $X2=0 $Y2=0
cc_203 N_A_284_21#_c_203_n N_A_27_47#_c_537_n 6.10702e-19 $X=1.995 $Y=1.185
+ $X2=0 $Y2=0
cc_204 N_A_284_21#_c_200_n N_A_27_47#_c_528_n 0.0114487f $X=1.495 $Y=1.185 $X2=0
+ $Y2=0
cc_205 N_A_284_21#_c_201_n N_A_27_47#_c_528_n 0.00370588f $X=1.92 $Y=1.26 $X2=0
+ $Y2=0
cc_206 N_A_284_21#_c_203_n N_A_27_47#_c_528_n 0.0129196f $X=1.995 $Y=1.185 $X2=0
+ $Y2=0
cc_207 N_A_284_21#_c_204_n N_A_27_47#_c_528_n 0.00492015f $X=2.605 $Y=1.26 $X2=0
+ $Y2=0
cc_208 N_A_284_21#_c_205_n N_A_27_47#_c_528_n 0.00161195f $X=2.68 $Y=1.185 $X2=0
+ $Y2=0
cc_209 N_A_284_21#_c_210_n N_A_27_47#_c_528_n 0.0102284f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_210 N_A_284_21#_c_200_n N_A_27_47#_c_529_n 0.00132005f $X=1.495 $Y=1.185
+ $X2=0 $Y2=0
cc_211 N_A_284_21#_c_200_n N_A_27_47#_c_530_n 6.46366e-19 $X=1.495 $Y=1.185
+ $X2=0 $Y2=0
cc_212 N_A_284_21#_c_203_n N_A_27_47#_c_530_n 0.0106336f $X=1.995 $Y=1.185 $X2=0
+ $Y2=0
cc_213 N_A_284_21#_c_228_p N_A_27_47#_c_530_n 0.0208586f $X=2.927 $Y=0.863 $X2=0
+ $Y2=0
cc_214 N_A_284_21#_c_208_n N_A_27_47#_c_530_n 0.0217594f $X=2.77 $Y=0.42 $X2=0
+ $Y2=0
cc_215 N_A_284_21#_c_209_n N_A_27_47#_c_530_n 0.00627978f $X=2.77 $Y=0.42 $X2=0
+ $Y2=0
cc_216 N_A_284_21#_c_200_n N_VGND_c_575_n 0.00373887f $X=1.495 $Y=1.185 $X2=0
+ $Y2=0
cc_217 N_A_284_21#_c_203_n N_VGND_c_575_n 0.00584655f $X=1.995 $Y=1.185 $X2=0
+ $Y2=0
cc_218 N_A_284_21#_c_208_n N_VGND_c_576_n 0.0561956f $X=2.77 $Y=0.42 $X2=0 $Y2=0
cc_219 N_A_284_21#_c_209_n N_VGND_c_576_n 0.00128418f $X=2.77 $Y=0.42 $X2=0
+ $Y2=0
cc_220 N_A_284_21#_c_200_n N_VGND_c_577_n 0.00547432f $X=1.495 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A_284_21#_c_203_n N_VGND_c_578_n 0.0054895f $X=1.995 $Y=1.185 $X2=0
+ $Y2=0
cc_222 N_A_284_21#_c_208_n N_VGND_c_578_n 0.0411871f $X=2.77 $Y=0.42 $X2=0 $Y2=0
cc_223 N_A_284_21#_c_209_n N_VGND_c_578_n 0.00215228f $X=2.77 $Y=0.42 $X2=0
+ $Y2=0
cc_224 N_A_284_21#_c_200_n N_VGND_c_580_n 0.0102326f $X=1.495 $Y=1.185 $X2=0
+ $Y2=0
cc_225 N_A_284_21#_c_203_n N_VGND_c_580_n 0.011357f $X=1.995 $Y=1.185 $X2=0
+ $Y2=0
cc_226 N_A_284_21#_c_208_n N_VGND_c_580_n 0.0228265f $X=2.77 $Y=0.42 $X2=0 $Y2=0
cc_227 N_TE_B_M1006_g N_A_M1011_g 0.0172168f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_228 N_TE_B_c_273_n N_A_M1011_g 4.68039e-19 $X=3.16 $Y=1.47 $X2=0 $Y2=0
cc_229 N_TE_B_M1008_g N_A_M1005_g 0.0167532f $X=3.25 $Y=0.905 $X2=0 $Y2=0
cc_230 N_TE_B_c_272_n N_A_c_351_n 0.0357822f $X=3.16 $Y=1.47 $X2=0 $Y2=0
cc_231 N_TE_B_c_273_n N_A_c_351_n 7.57433e-19 $X=3.16 $Y=1.47 $X2=0 $Y2=0
cc_232 N_TE_B_M1006_g N_A_c_352_n 5.06247e-19 $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_233 N_TE_B_c_272_n N_A_c_352_n 0.00422393f $X=3.16 $Y=1.47 $X2=0 $Y2=0
cc_234 N_TE_B_c_273_n N_A_c_352_n 0.0656317f $X=3.16 $Y=1.47 $X2=0 $Y2=0
cc_235 N_TE_B_c_274_n N_A_39_367#_c_387_n 9.91822e-19 $X=1.415 $Y=1.725 $X2=0
+ $Y2=0
cc_236 N_TE_B_c_274_n N_A_39_367#_c_398_n 0.0144236f $X=1.415 $Y=1.725 $X2=0
+ $Y2=0
cc_237 N_TE_B_c_277_n N_A_39_367#_c_398_n 6.58365e-19 $X=1.845 $Y=1.725 $X2=0
+ $Y2=0
cc_238 N_TE_B_c_274_n N_A_39_367#_c_388_n 0.0111508f $X=1.415 $Y=1.725 $X2=0
+ $Y2=0
cc_239 N_TE_B_c_267_n N_A_39_367#_c_388_n 0.00212913f $X=1.77 $Y=1.65 $X2=0
+ $Y2=0
cc_240 N_TE_B_c_277_n N_A_39_367#_c_388_n 0.0111561f $X=1.845 $Y=1.725 $X2=0
+ $Y2=0
cc_241 N_TE_B_c_277_n N_A_39_367#_c_389_n 0.00110817f $X=1.845 $Y=1.725 $X2=0
+ $Y2=0
cc_242 N_TE_B_c_269_n N_A_39_367#_c_389_n 0.0030275f $X=2.995 $Y=1.65 $X2=0
+ $Y2=0
cc_243 N_TE_B_c_274_n N_A_39_367#_c_403_n 7.12253e-19 $X=1.415 $Y=1.725 $X2=0
+ $Y2=0
cc_244 N_TE_B_c_277_n N_A_39_367#_c_403_n 0.0154933f $X=1.845 $Y=1.725 $X2=0
+ $Y2=0
cc_245 N_TE_B_c_273_n N_VPWR_M1006_d 0.00188947f $X=3.16 $Y=1.47 $X2=0 $Y2=0
cc_246 N_TE_B_c_274_n N_VPWR_c_473_n 0.00372815f $X=1.415 $Y=1.725 $X2=0 $Y2=0
cc_247 N_TE_B_c_277_n N_VPWR_c_473_n 0.00372815f $X=1.845 $Y=1.725 $X2=0 $Y2=0
cc_248 N_TE_B_M1006_g N_VPWR_c_474_n 0.00307315f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_249 N_TE_B_c_277_n N_VPWR_c_475_n 0.0054895f $X=1.845 $Y=1.725 $X2=0 $Y2=0
cc_250 N_TE_B_M1006_g N_VPWR_c_475_n 0.00343766f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_251 N_TE_B_c_274_n N_VPWR_c_477_n 0.00547432f $X=1.415 $Y=1.725 $X2=0 $Y2=0
cc_252 N_TE_B_c_274_n N_VPWR_c_472_n 0.00978129f $X=1.415 $Y=1.725 $X2=0 $Y2=0
cc_253 N_TE_B_c_277_n N_VPWR_c_472_n 0.0110927f $X=1.845 $Y=1.725 $X2=0 $Y2=0
cc_254 N_TE_B_M1006_g N_VPWR_c_472_n 0.00489211f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_255 N_TE_B_c_267_n N_A_27_47#_c_528_n 3.53029e-19 $X=1.77 $Y=1.65 $X2=0 $Y2=0
cc_256 N_TE_B_c_269_n N_A_27_47#_c_528_n 3.5987e-19 $X=2.995 $Y=1.65 $X2=0 $Y2=0
cc_257 N_TE_B_c_268_n N_A_27_47#_c_529_n 3.55022e-19 $X=1.49 $Y=1.65 $X2=0 $Y2=0
cc_258 N_TE_B_M1008_g N_VGND_c_576_n 0.00395118f $X=3.25 $Y=0.905 $X2=0 $Y2=0
cc_259 N_TE_B_M1008_g N_VGND_c_578_n 0.00326842f $X=3.25 $Y=0.905 $X2=0 $Y2=0
cc_260 N_TE_B_M1008_g N_VGND_c_580_n 0.00378428f $X=3.25 $Y=0.905 $X2=0 $Y2=0
cc_261 N_A_M1011_g N_VPWR_c_474_n 0.00924062f $X=3.785 $Y=2.775 $X2=0 $Y2=0
cc_262 N_A_M1011_g N_VPWR_c_478_n 0.00424868f $X=3.785 $Y=2.775 $X2=0 $Y2=0
cc_263 N_A_M1011_g N_VPWR_c_472_n 0.00839126f $X=3.785 $Y=2.775 $X2=0 $Y2=0
cc_264 N_A_M1005_g N_VGND_c_576_n 0.00613414f $X=3.82 $Y=0.905 $X2=0 $Y2=0
cc_265 N_A_c_351_n N_VGND_c_576_n 0.00104907f $X=3.73 $Y=1.47 $X2=0 $Y2=0
cc_266 N_A_c_352_n N_VGND_c_576_n 0.0174749f $X=3.73 $Y=1.47 $X2=0 $Y2=0
cc_267 N_A_M1005_g N_VGND_c_579_n 0.00366993f $X=3.82 $Y=0.905 $X2=0 $Y2=0
cc_268 N_A_M1005_g N_VGND_c_580_n 0.0045051f $X=3.82 $Y=0.905 $X2=0 $Y2=0
cc_269 N_A_39_367#_c_393_n N_Z_M1002_d 0.00332344f $X=1.035 $Y=2.99 $X2=0 $Y2=0
cc_270 N_A_39_367#_M1002_s N_Z_c_440_n 7.12223e-19 $X=0.195 $Y=1.835 $X2=0 $Y2=0
cc_271 N_A_39_367#_c_386_n N_Z_c_440_n 0.00728199f $X=0.34 $Y=2.22 $X2=0 $Y2=0
cc_272 N_A_39_367#_c_387_n N_Z_c_440_n 0.00691492f $X=1.2 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_39_367#_M1002_s N_Z_c_441_n 0.00252613f $X=0.195 $Y=1.835 $X2=0 $Y2=0
cc_274 N_A_39_367#_c_386_n N_Z_c_441_n 0.0162061f $X=0.34 $Y=2.22 $X2=0 $Y2=0
cc_275 N_A_39_367#_c_393_n N_Z_c_461_n 0.0126348f $X=1.035 $Y=2.99 $X2=0 $Y2=0
cc_276 N_A_39_367#_c_388_n N_VPWR_M1000_s 0.00176461f $X=1.895 $Y=1.9 $X2=-0.19
+ $Y2=1.655
cc_277 N_A_39_367#_c_388_n N_VPWR_c_473_n 0.0135055f $X=1.895 $Y=1.9 $X2=0 $Y2=0
cc_278 N_A_39_367#_c_403_n N_VPWR_c_475_n 0.0153681f $X=2.06 $Y=2.91 $X2=0 $Y2=0
cc_279 N_A_39_367#_c_385_n N_VPWR_c_477_n 0.021159f $X=0.34 $Y=2.905 $X2=0 $Y2=0
cc_280 N_A_39_367#_c_393_n N_VPWR_c_477_n 0.0298674f $X=1.035 $Y=2.99 $X2=0
+ $Y2=0
cc_281 N_A_39_367#_c_398_n N_VPWR_c_477_n 0.01906f $X=1.2 $Y=2.905 $X2=0 $Y2=0
cc_282 N_A_39_367#_M1002_s N_VPWR_c_472_n 0.00231914f $X=0.195 $Y=1.835 $X2=0
+ $Y2=0
cc_283 N_A_39_367#_M1010_s N_VPWR_c_472_n 0.00223559f $X=1.06 $Y=1.835 $X2=0
+ $Y2=0
cc_284 N_A_39_367#_M1003_d N_VPWR_c_472_n 0.00444118f $X=1.92 $Y=1.835 $X2=0
+ $Y2=0
cc_285 N_A_39_367#_c_385_n N_VPWR_c_472_n 0.0126421f $X=0.34 $Y=2.905 $X2=0
+ $Y2=0
cc_286 N_A_39_367#_c_393_n N_VPWR_c_472_n 0.0187823f $X=1.035 $Y=2.99 $X2=0
+ $Y2=0
cc_287 N_A_39_367#_c_398_n N_VPWR_c_472_n 0.0124545f $X=1.2 $Y=2.905 $X2=0 $Y2=0
cc_288 N_A_39_367#_c_403_n N_VPWR_c_472_n 0.00945867f $X=2.06 $Y=2.91 $X2=0
+ $Y2=0
cc_289 N_Z_M1002_d N_VPWR_c_472_n 0.00225186f $X=0.63 $Y=1.835 $X2=0 $Y2=0
cc_290 N_Z_c_437_n N_A_27_47#_M1001_s 7.12223e-19 $X=0.615 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_291 N_Z_c_438_n N_A_27_47#_M1001_s 0.00353051f $X=0.355 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_292 N_Z_c_437_n N_A_27_47#_c_526_n 0.00538516f $X=0.615 $Y=1.04 $X2=0 $Y2=0
cc_293 N_Z_c_438_n N_A_27_47#_c_526_n 0.0203954f $X=0.355 $Y=1.04 $X2=0 $Y2=0
cc_294 N_Z_M1001_d N_A_27_47#_c_531_n 0.00352365f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_295 N_Z_c_437_n N_A_27_47#_c_531_n 0.00359356f $X=0.615 $Y=1.04 $X2=0 $Y2=0
cc_296 N_Z_c_451_n N_A_27_47#_c_531_n 0.0157977f $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_297 N_Z_c_437_n N_A_27_47#_c_529_n 0.00948931f $X=0.615 $Y=1.04 $X2=0 $Y2=0
cc_298 N_Z_M1001_d N_VGND_c_580_n 0.00233228f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_299 N_A_27_47#_c_528_n N_VGND_M1004_s 0.00250873f $X=2.045 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_300 N_A_27_47#_c_528_n N_VGND_c_575_n 0.0192006f $X=2.045 $Y=1.04 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_531_n N_VGND_c_577_n 0.0364508f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_527_n N_VGND_c_577_n 0.022075f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_536_n N_VGND_c_577_n 0.0207136f $X=1.28 $Y=0.425 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_530_n N_VGND_c_578_n 0.0210192f $X=2.21 $Y=0.42 $X2=0 $Y2=0
cc_305 N_A_27_47#_M1001_s N_VGND_c_580_n 0.00282988f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1009_s N_VGND_c_580_n 0.00280658f $X=1.07 $Y=0.235 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_M1007_d N_VGND_c_580_n 0.00231914f $X=2.07 $Y=0.235 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_531_n N_VGND_c_580_n 0.0238173f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_309 N_A_27_47#_c_527_n N_VGND_c_580_n 0.0127477f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_536_n N_VGND_c_580_n 0.0126421f $X=1.28 $Y=0.425 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_530_n N_VGND_c_580_n 0.0125689f $X=2.21 $Y=0.42 $X2=0 $Y2=0
