* File: sky130_fd_sc_lp__o41ai_0.spice
* Created: Fri Aug 28 11:20:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o41ai_0  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_A_218_57#_M1006_d N_B1_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.3087 PD=0.7 PS=2.31 NRD=0 NRS=194.28 M=1 R=2.8 SA=75000.7
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A4_M1001_g N_A_218_57#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07875 AS=0.0588 PD=0.795 PS=0.7 NRD=12.852 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_218_57#_M1002_d N_A3_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.07875 PD=0.7 PS=0.795 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_218_57#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0588 PD=0.755 PS=0.7 NRD=8.568 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_218_57#_M1005_d N_A1_M1005_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.07035 PD=1.37 PS=0.755 NRD=0 NRS=7.14 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1004 A_291_483# N_A4_M1004_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=0.64 AD=0.1168
+ AS=0.0896 PD=1.005 PS=0.92 NRD=39.2424 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1003 A_394_483# N_A3_M1003_g A_291_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.096
+ AS=0.1168 PD=0.94 PS=1.005 NRD=29.2348 NRS=39.2424 M=1 R=4.26667 SA=75001.1
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1007 A_484_483# N_A2_M1007_g A_394_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.096 PD=0.85 PS=0.94 NRD=15.3857 NRS=29.2348 M=1 R=4.26667 SA=75001.6
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_484_483# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_77 VPB 0 9.44548e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o41ai_0.pxi.spice"
*
.ends
*
*
