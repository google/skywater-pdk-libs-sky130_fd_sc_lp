* File: sky130_fd_sc_lp__dlxtn_1.spice
* Created: Wed Sep  2 09:48:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxtn_1.pex.spice"
.subckt sky130_fd_sc_lp__dlxtn_1  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_D_M1009_g N_A_59_129#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_228_129#_M1004_d N_GATE_N_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_228_129#_M1011_g N_A_342_481#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1003 A_656_47# N_A_59_129#_M1003_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1016 N_A_656_481#_M1016_d N_A_228_129#_M1016_g A_656_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1008 A_836_47# N_A_342_481#_M1008_g N_A_656_481#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_842_413#_M1014_g A_836_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.0819 PD=0.81 PS=0.81 NRD=18.564 NRS=39.996 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_842_413#_M1017_d N_A_656_481#_M1017_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=2.136 M=1 R=5.6
+ SA=75001.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_Q_M1006_d N_A_842_413#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_D_M1001_g N_A_59_129#_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_A_228_129#_M1005_d N_GATE_N_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_228_129#_M1000_g N_A_342_481#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2064 AS=0.1696 PD=1.285 PS=1.81 NRD=83.0946 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1012 A_584_481# N_A_59_129#_M1012_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.2064 PD=0.85 PS=1.285 NRD=15.3857 NRS=29.2348 M=1 R=4.26667
+ SA=75001 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1013 N_A_656_481#_M1013_d N_A_342_481#_M1013_g A_584_481# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1002 A_764_481# N_A_228_129#_M1002_g N_A_656_481#_M1013_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0880019 PD=0.81 PS=0.816226 NRD=65.6601 NRS=53.9386 M=1
+ R=2.8 SA=75001.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_842_413#_M1007_g A_764_481# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.144375 AS=0.0819 PD=1.0525 PS=0.81 NRD=267.349 NRS=65.6601 M=1 R=2.8
+ SA=75002.4 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_842_413#_M1010_d N_A_656_481#_M1010_g N_VPWR_M1007_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.433125 PD=3.05 PS=3.1575 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.3 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1015 N_Q_M1015_d N_A_842_413#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=13.3351 P=18.11
*
.include "sky130_fd_sc_lp__dlxtn_1.pxi.spice"
*
.ends
*
*
