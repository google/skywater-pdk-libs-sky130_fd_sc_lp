# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.925000 1.315000 1.045000 ;
        RECT 1.065000 1.045000 2.245000 1.790000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.365000 1.605000 8.505000 1.775000 ;
        RECT 7.365000 1.775000 7.610000 3.075000 ;
        RECT 7.445000 0.255000 7.635000 0.845000 ;
        RECT 7.445000 0.845000 8.505000 1.015000 ;
        RECT 8.210000 1.775000 8.505000 2.470000 ;
        RECT 8.210000 2.470000 8.445000 3.075000 ;
        RECT 8.305000 0.425000 8.505000 0.845000 ;
        RECT 8.305000 1.015000 8.505000 1.605000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.435000 2.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.474000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.210000 6.085000 1.760000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  2.660000 0.365000 3.245000 ;
      RECT 0.205000  0.085000 0.535000 0.670000 ;
      RECT 0.705000  0.395000 0.975000 0.725000 ;
      RECT 0.705000  0.725000 0.895000 1.960000 ;
      RECT 0.705000  1.960000 2.045000 2.130000 ;
      RECT 0.705000  2.130000 1.215000 2.990000 ;
      RECT 1.170000  0.085000 1.480000 0.725000 ;
      RECT 1.445000  2.300000 1.705000 3.245000 ;
      RECT 1.650000  0.395000 1.980000 0.615000 ;
      RECT 1.650000  0.615000 2.605000 0.785000 ;
      RECT 1.875000  2.130000 2.045000 2.885000 ;
      RECT 1.875000  2.885000 3.010000 3.075000 ;
      RECT 2.225000  2.045000 2.605000 2.715000 ;
      RECT 2.265000  0.255000 3.870000 0.445000 ;
      RECT 2.425000  0.785000 2.605000 2.045000 ;
      RECT 2.775000  0.710000 3.010000 2.885000 ;
      RECT 3.180000  0.710000 3.475000 1.250000 ;
      RECT 3.180000  1.250000 4.540000 1.465000 ;
      RECT 3.180000  1.465000 3.475000 2.695000 ;
      RECT 3.700000  0.445000 3.870000 0.525000 ;
      RECT 3.700000  0.525000 5.430000 0.695000 ;
      RECT 3.805000  1.635000 4.915000 1.805000 ;
      RECT 3.805000  1.805000 4.140000 2.095000 ;
      RECT 3.935000  2.360000 4.530000 3.245000 ;
      RECT 4.050000  0.085000 4.380000 0.355000 ;
      RECT 4.340000  1.985000 4.530000 2.360000 ;
      RECT 4.560000  0.865000 4.915000 1.080000 ;
      RECT 4.710000  1.805000 4.915000 2.310000 ;
      RECT 4.710000  2.310000 6.075000 2.490000 ;
      RECT 4.710000  2.490000 5.040000 2.930000 ;
      RECT 4.720000  1.080000 4.915000 1.635000 ;
      RECT 5.085000  0.270000 5.430000 0.525000 ;
      RECT 5.085000  0.695000 5.255000 1.930000 ;
      RECT 5.085000  1.930000 5.725000 2.140000 ;
      RECT 5.625000  0.085000 5.955000 1.040000 ;
      RECT 5.905000  1.930000 6.435000 2.100000 ;
      RECT 5.905000  2.100000 6.075000 2.310000 ;
      RECT 5.980000  2.785000 6.190000 3.245000 ;
      RECT 6.265000  1.345000 6.855000 1.675000 ;
      RECT 6.265000  1.675000 6.435000 1.930000 ;
      RECT 6.410000  2.280000 6.785000 2.950000 ;
      RECT 6.415000  0.255000 6.685000 0.995000 ;
      RECT 6.415000  0.995000 7.195000 1.175000 ;
      RECT 6.615000  1.845000 7.195000 2.015000 ;
      RECT 6.615000  2.015000 6.785000 2.280000 ;
      RECT 6.945000  0.085000 7.275000 0.825000 ;
      RECT 6.955000  2.185000 7.195000 3.245000 ;
      RECT 7.025000  1.175000 7.195000 1.185000 ;
      RECT 7.025000  1.185000 8.135000 1.435000 ;
      RECT 7.025000  1.435000 7.195000 1.845000 ;
      RECT 7.780000  1.945000 8.040000 3.245000 ;
      RECT 7.805000  0.085000 8.135000 0.675000 ;
      RECT 8.675000  0.085000 8.995000 1.090000 ;
      RECT 8.675000  1.815000 8.935000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__sdlclkp_4
END LIBRARY
