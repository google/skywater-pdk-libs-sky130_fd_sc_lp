* File: sky130_fd_sc_lp__ha_1.spice
* Created: Wed Sep  2 09:54:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ha_1.pex.spice"
.subckt sky130_fd_sc_lp__ha_1  VNB VPB B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_80_30#_M1009_g N_SUM_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_307_62#_M1007_d N_A_223_320#_M1007_g N_A_80_30#_M1007_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_B_M1012_g N_A_307_62#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_307_62#_M1004_d N_A_M1004_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1010 A_675_146# N_B_M1010_g N_A_223_320#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g A_675_146# VNB NSHORT L=0.15 W=0.42 AD=0.0896
+ AS=0.0504 PD=0.81 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1013 N_COUT_M1013_d N_A_223_320#_M1013_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=3.204 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_30#_M1003_g N_SUM_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.398475 AS=0.3339 PD=2.9925 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1008 N_A_80_30#_M1008_d N_A_223_320#_M1008_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.132825 PD=0.7 PS=0.9975 NRD=0 NRS=215.754 M=1 R=2.8
+ SA=75001.1 SB=75003 A=0.063 P=1.14 MULT=1
MM1002 A_401_428# N_B_M1002_g N_A_80_30#_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0588 PD=0.8 PS=0.7 NRD=63.3158 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g A_401_428# VPB PHIGHVT L=0.15 W=0.42 AD=0.1449
+ AS=0.0798 PD=1.11 PS=0.8 NRD=23.443 NRS=63.3158 M=1 R=2.8 SA=75002 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_223_320#_M1006_d N_B_M1006_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1449 PD=0.7 PS=1.11 NRD=0 NRS=0 M=1 R=2.8 SA=75002.9 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_223_320#_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.099225 AS=0.0588 PD=0.8375 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.3
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_COUT_M1001_d N_A_223_320#_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.297675 PD=3.05 PS=2.5125 NRD=0 NRS=7.0329 M=1 R=8.4
+ SA=75001.4 SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__ha_1.pxi.spice"
*
.ends
*
*
