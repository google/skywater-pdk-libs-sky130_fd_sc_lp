* File: sky130_fd_sc_lp__o41ai_lp.pxi.spice
* Created: Fri Aug 28 11:20:43 2020
* 
x_PM_SKY130_FD_SC_LP__O41AI_LP%B1 N_B1_M1002_g N_B1_M1007_g N_B1_c_67_n
+ N_B1_c_68_n B1 B1 N_B1_c_69_n N_B1_c_70_n PM_SKY130_FD_SC_LP__O41AI_LP%B1
x_PM_SKY130_FD_SC_LP__O41AI_LP%A4 N_A4_M1003_g N_A4_c_103_n N_A4_M1009_g
+ N_A4_c_104_n A4 A4 N_A4_c_106_n PM_SKY130_FD_SC_LP__O41AI_LP%A4
x_PM_SKY130_FD_SC_LP__O41AI_LP%A3 N_A3_M1001_g N_A3_M1000_g N_A3_c_149_n
+ N_A3_c_154_n A3 A3 A3 A3 N_A3_c_150_n N_A3_c_151_n
+ PM_SKY130_FD_SC_LP__O41AI_LP%A3
x_PM_SKY130_FD_SC_LP__O41AI_LP%A2 N_A2_M1004_g N_A2_M1008_g N_A2_c_198_n
+ N_A2_c_203_n A2 A2 A2 A2 N_A2_c_199_n N_A2_c_200_n
+ PM_SKY130_FD_SC_LP__O41AI_LP%A2
x_PM_SKY130_FD_SC_LP__O41AI_LP%A1 N_A1_M1006_g N_A1_M1005_g A1 N_A1_c_244_n
+ PM_SKY130_FD_SC_LP__O41AI_LP%A1
x_PM_SKY130_FD_SC_LP__O41AI_LP%VPWR N_VPWR_M1002_s N_VPWR_M1006_d N_VPWR_c_272_n
+ N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n VPWR N_VPWR_c_276_n
+ N_VPWR_c_271_n PM_SKY130_FD_SC_LP__O41AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O41AI_LP%Y N_Y_M1007_s N_Y_M1002_d N_Y_c_310_n N_Y_c_313_n
+ N_Y_c_314_n N_Y_c_322_n Y N_Y_c_311_n PM_SKY130_FD_SC_LP__O41AI_LP%Y
x_PM_SKY130_FD_SC_LP__O41AI_LP%A_153_57# N_A_153_57#_M1007_d N_A_153_57#_M1000_d
+ N_A_153_57#_M1005_d N_A_153_57#_c_353_n N_A_153_57#_c_354_n
+ N_A_153_57#_c_355_n N_A_153_57#_c_356_n N_A_153_57#_c_357_n
+ N_A_153_57#_c_358_n N_A_153_57#_c_359_n PM_SKY130_FD_SC_LP__O41AI_LP%A_153_57#
x_PM_SKY130_FD_SC_LP__O41AI_LP%VGND N_VGND_M1003_d N_VGND_M1004_d N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ VGND N_VGND_c_416_n N_VGND_c_417_n PM_SKY130_FD_SC_LP__O41AI_LP%VGND
cc_1 VNB N_B1_M1007_g 0.0370962f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.495
cc_2 VNB N_B1_c_67_n 0.0234927f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.63
cc_3 VNB N_B1_c_68_n 0.00173762f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.795
cc_4 VNB N_B1_c_69_n 0.0165772f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_5 VNB N_B1_c_70_n 0.00737816f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_6 VNB N_A4_M1003_g 0.0350627f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.595
cc_7 VNB N_A4_c_103_n 0.00170515f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.125
cc_8 VNB N_A4_c_104_n 0.0230536f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.63
cc_9 VNB A4 0.0017033f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.795
cc_10 VNB N_A4_c_106_n 0.0171231f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_11 VNB N_A3_M1000_g 0.0424525f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.495
cc_12 VNB N_A3_c_149_n 0.0155516f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.63
cc_13 VNB N_A3_c_150_n 0.0165355f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.295
cc_14 VNB N_A3_c_151_n 0.00207575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_M1004_g 0.0420602f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.595
cc_16 VNB N_A2_c_198_n 0.0144577f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.63
cc_17 VNB N_A2_c_199_n 0.0157585f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.295
cc_18 VNB N_A2_c_200_n 0.00488064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1005_g 0.0525284f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.495
cc_20 VNB A1 0.0197399f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_21 VNB N_A1_c_244_n 0.0490242f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.795
cc_22 VNB N_VPWR_c_271_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_310_n 0.0449558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_311_n 0.0319193f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_25 VNB N_A_153_57#_c_353_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.795
cc_26 VNB N_A_153_57#_c_354_n 0.0155653f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB N_A_153_57#_c_355_n 0.00812185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_153_57#_c_356_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_29 VNB N_A_153_57#_c_357_n 0.0267662f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.29
cc_30 VNB N_A_153_57#_c_358_n 0.0261109f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.665
cc_31 VNB N_A_153_57#_c_359_n 0.00828526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_410_n 0.00714888f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_33 VNB N_VGND_c_411_n 0.00712794f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_34 VNB N_VGND_c_412_n 0.0348078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_413_n 0.00632158f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_36 VNB N_VGND_c_414_n 0.0204586f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_37 VNB N_VGND_c_415_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.29
cc_38 VNB N_VGND_c_416_n 0.0217109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_417_n 0.211282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_B1_M1002_g 0.0379906f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.595
cc_41 VPB N_B1_c_68_n 0.0119856f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.795
cc_42 VPB N_B1_c_70_n 0.00190365f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.29
cc_43 VPB N_A4_c_103_n 0.0117752f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.125
cc_44 VPB N_A4_M1009_g 0.0338012f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.495
cc_45 VPB A4 0.00195814f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.795
cc_46 VPB N_A3_M1001_g 0.0250137f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.595
cc_47 VPB N_A3_c_149_n 0.00791466f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.63
cc_48 VPB N_A3_c_154_n 0.0139631f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.795
cc_49 VPB N_A3_c_151_n 0.00102431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A2_M1008_g 0.0248471f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.495
cc_51 VPB N_A2_c_198_n 0.00735792f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.63
cc_52 VPB N_A2_c_203_n 0.0129076f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.795
cc_53 VPB N_A2_c_200_n 0.00453314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A1_M1006_g 0.0361751f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.595
cc_55 VPB A1 0.010102f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.29
cc_56 VPB N_A1_c_244_n 0.0280935f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.795
cc_57 VPB N_VPWR_c_272_n 0.0140081f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.495
cc_58 VPB N_VPWR_c_273_n 0.0320215f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.29
cc_59 VPB N_VPWR_c_274_n 0.0110854f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.63
cc_60 VPB N_VPWR_c_275_n 0.0436066f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_61 VPB N_VPWR_c_276_n 0.0655349f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.29
cc_62 VPB N_VPWR_c_271_n 0.0492815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_Y_c_310_n 0.0155974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_Y_c_313_n 0.0148215f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.29
cc_65 VPB N_Y_c_314_n 0.0119416f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.125
cc_66 N_B1_M1007_g N_A4_M1003_g 0.0276106f $X=0.69 $Y=0.495 $X2=0 $Y2=0
cc_67 N_B1_c_68_n N_A4_c_103_n 0.0139409f $X=0.63 $Y=1.795 $X2=0 $Y2=0
cc_68 N_B1_M1002_g N_A4_M1009_g 0.0341185f $X=0.64 $Y=2.595 $X2=0 $Y2=0
cc_69 N_B1_c_67_n N_A4_c_104_n 0.0139409f $X=0.63 $Y=1.63 $X2=0 $Y2=0
cc_70 N_B1_c_69_n A4 7.89554e-19 $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_71 N_B1_c_70_n A4 0.0510782f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_72 N_B1_c_69_n N_A4_c_106_n 0.0139409f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_73 N_B1_c_70_n N_A4_c_106_n 0.00382187f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_74 N_B1_M1002_g N_VPWR_c_273_n 0.0208226f $X=0.64 $Y=2.595 $X2=0 $Y2=0
cc_75 N_B1_M1002_g N_VPWR_c_276_n 0.00840199f $X=0.64 $Y=2.595 $X2=0 $Y2=0
cc_76 N_B1_M1002_g N_VPWR_c_271_n 0.0136033f $X=0.64 $Y=2.595 $X2=0 $Y2=0
cc_77 N_B1_M1002_g N_Y_c_310_n 0.00609602f $X=0.64 $Y=2.595 $X2=0 $Y2=0
cc_78 N_B1_M1007_g N_Y_c_310_n 0.0091713f $X=0.69 $Y=0.495 $X2=0 $Y2=0
cc_79 N_B1_c_69_n N_Y_c_310_n 0.0148853f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_80 N_B1_c_70_n N_Y_c_310_n 0.0484816f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_81 N_B1_M1002_g N_Y_c_313_n 0.0216533f $X=0.64 $Y=2.595 $X2=0 $Y2=0
cc_82 N_B1_c_68_n N_Y_c_313_n 5.70285e-19 $X=0.63 $Y=1.795 $X2=0 $Y2=0
cc_83 N_B1_c_70_n N_Y_c_313_n 0.0272409f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_84 N_B1_M1002_g N_Y_c_322_n 0.0243371f $X=0.64 $Y=2.595 $X2=0 $Y2=0
cc_85 N_B1_M1007_g N_Y_c_311_n 0.0089501f $X=0.69 $Y=0.495 $X2=0 $Y2=0
cc_86 N_B1_c_69_n N_Y_c_311_n 6.1174e-19 $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_87 N_B1_c_70_n N_Y_c_311_n 0.00422224f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_88 N_B1_M1007_g N_A_153_57#_c_353_n 0.00747924f $X=0.69 $Y=0.495 $X2=0 $Y2=0
cc_89 N_B1_M1007_g N_A_153_57#_c_355_n 0.00539129f $X=0.69 $Y=0.495 $X2=0 $Y2=0
cc_90 N_B1_c_69_n N_A_153_57#_c_355_n 2.31969e-19 $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_91 N_B1_c_70_n N_A_153_57#_c_355_n 0.00718195f $X=0.63 $Y=1.29 $X2=0 $Y2=0
cc_92 N_B1_M1007_g N_VGND_c_412_n 0.00502664f $X=0.69 $Y=0.495 $X2=0 $Y2=0
cc_93 N_B1_M1007_g N_VGND_c_417_n 0.0103055f $X=0.69 $Y=0.495 $X2=0 $Y2=0
cc_94 N_A4_M1003_g N_A3_M1000_g 0.0197176f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_95 A4 N_A3_M1000_g 8.29967e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A4_c_106_n N_A3_M1000_g 0.00528503f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_97 N_A4_c_104_n N_A3_c_149_n 0.0107256f $X=1.17 $Y=1.63 $X2=0 $Y2=0
cc_98 N_A4_c_103_n N_A3_c_154_n 0.0107256f $X=1.17 $Y=1.795 $X2=0 $Y2=0
cc_99 N_A4_M1009_g N_A3_c_154_n 0.0744221f $X=1.17 $Y=2.595 $X2=0 $Y2=0
cc_100 A4 N_A3_c_150_n 0.00183897f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A4_c_106_n N_A3_c_150_n 0.0107256f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_102 N_A4_M1009_g N_A3_c_151_n 0.00489631f $X=1.17 $Y=2.595 $X2=0 $Y2=0
cc_103 A4 N_A3_c_151_n 0.0334612f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A4_c_106_n N_A3_c_151_n 0.00183897f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_105 N_A4_M1009_g N_VPWR_c_273_n 0.00121833f $X=1.17 $Y=2.595 $X2=0 $Y2=0
cc_106 N_A4_M1009_g N_VPWR_c_276_n 0.00939541f $X=1.17 $Y=2.595 $X2=0 $Y2=0
cc_107 N_A4_M1009_g N_VPWR_c_271_n 0.0161801f $X=1.17 $Y=2.595 $X2=0 $Y2=0
cc_108 N_A4_c_103_n N_Y_c_313_n 3.03142e-19 $X=1.17 $Y=1.795 $X2=0 $Y2=0
cc_109 N_A4_M1009_g N_Y_c_313_n 0.00498701f $X=1.17 $Y=2.595 $X2=0 $Y2=0
cc_110 A4 N_Y_c_313_n 0.00534367f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A4_M1009_g N_Y_c_322_n 0.0208563f $X=1.17 $Y=2.595 $X2=0 $Y2=0
cc_112 N_A4_M1003_g N_A_153_57#_c_353_n 0.00893067f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_113 N_A4_M1003_g N_A_153_57#_c_354_n 0.00933704f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_114 A4 N_A_153_57#_c_354_n 0.019672f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A4_c_106_n N_A_153_57#_c_354_n 9.55426e-19 $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_116 N_A4_M1003_g N_A_153_57#_c_355_n 0.0027409f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_117 A4 N_A_153_57#_c_355_n 0.00534367f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_A4_c_106_n N_A_153_57#_c_355_n 3.01559e-19 $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_119 N_A4_M1003_g N_A_153_57#_c_356_n 8.62854e-19 $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_120 N_A4_M1003_g N_A_153_57#_c_359_n 4.36217e-19 $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_121 N_A4_M1003_g N_VGND_c_410_n 0.00503903f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_122 N_A4_M1003_g N_VGND_c_412_n 0.00502664f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_123 N_A4_M1003_g N_VGND_c_417_n 0.00585942f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_124 N_A3_M1000_g N_A2_M1004_g 0.0340643f $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_125 N_A3_M1001_g N_A2_M1008_g 0.051978f $X=1.67 $Y=2.595 $X2=0 $Y2=0
cc_126 N_A3_c_151_n N_A2_M1008_g 0.00303803f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_127 N_A3_c_149_n N_A2_c_198_n 0.0117523f $X=1.71 $Y=1.77 $X2=0 $Y2=0
cc_128 N_A3_c_154_n N_A2_c_203_n 0.0117523f $X=1.71 $Y=1.935 $X2=0 $Y2=0
cc_129 N_A3_c_150_n N_A2_c_199_n 0.0117523f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_130 N_A3_c_151_n N_A2_c_199_n 7.56445e-19 $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_131 N_A3_M1001_g N_A2_c_200_n 0.0029856f $X=1.67 $Y=2.595 $X2=0 $Y2=0
cc_132 N_A3_c_150_n N_A2_c_200_n 0.00411743f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_133 N_A3_c_151_n N_A2_c_200_n 0.12625f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_134 N_A3_M1001_g N_VPWR_c_276_n 0.00656883f $X=1.67 $Y=2.595 $X2=0 $Y2=0
cc_135 N_A3_c_151_n N_VPWR_c_276_n 0.00914393f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_136 N_A3_M1001_g N_VPWR_c_271_n 0.00827299f $X=1.67 $Y=2.595 $X2=0 $Y2=0
cc_137 N_A3_c_151_n N_VPWR_c_271_n 0.0101955f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_138 N_A3_M1001_g N_Y_c_313_n 4.29532e-19 $X=1.67 $Y=2.595 $X2=0 $Y2=0
cc_139 N_A3_c_151_n N_Y_c_313_n 0.00586766f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_140 N_A3_M1001_g N_Y_c_322_n 0.00264353f $X=1.67 $Y=2.595 $X2=0 $Y2=0
cc_141 N_A3_c_151_n N_Y_c_322_n 0.0242282f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_142 N_A3_c_151_n A_359_419# 0.00742697f $X=1.71 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_143 N_A3_M1000_g N_A_153_57#_c_353_n 8.47653e-19 $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_144 N_A3_M1000_g N_A_153_57#_c_354_n 0.00998365f $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_145 N_A3_c_150_n N_A_153_57#_c_354_n 8.47771e-19 $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_146 N_A3_c_151_n N_A_153_57#_c_354_n 0.0126089f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_147 N_A3_M1000_g N_A_153_57#_c_356_n 0.00933335f $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_148 N_A3_M1000_g N_A_153_57#_c_359_n 0.00629384f $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_149 N_A3_c_150_n N_A_153_57#_c_359_n 2.96131e-19 $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_150 N_A3_c_151_n N_A_153_57#_c_359_n 0.00458006f $X=1.71 $Y=1.43 $X2=0 $Y2=0
cc_151 N_A3_M1000_g N_VGND_c_410_n 0.00579413f $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_152 N_A3_M1000_g N_VGND_c_414_n 0.00502664f $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_153 N_A3_M1000_g N_VGND_c_417_n 0.00597972f $X=1.76 $Y=0.495 $X2=0 $Y2=0
cc_154 N_A2_M1008_g N_A1_M1006_g 0.0488274f $X=2.24 $Y=2.595 $X2=0 $Y2=0
cc_155 N_A2_c_198_n N_A1_M1006_g 0.0182716f $X=2.28 $Y=1.77 $X2=0 $Y2=0
cc_156 N_A2_c_200_n N_A1_M1006_g 0.0108706f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_157 N_A2_M1004_g N_A1_M1005_g 0.02501f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_158 N_A2_c_199_n A1 0.00191036f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_159 N_A2_c_200_n A1 0.0264142f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_160 N_A2_M1004_g N_A1_c_244_n 0.00132528f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_161 N_A2_c_199_n N_A1_c_244_n 0.0182716f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_162 N_A2_c_200_n N_A1_c_244_n 0.00291303f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_163 N_A2_M1008_g N_VPWR_c_275_n 0.00238668f $X=2.24 $Y=2.595 $X2=0 $Y2=0
cc_164 N_A2_c_200_n N_VPWR_c_275_n 0.0294543f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_165 N_A2_M1008_g N_VPWR_c_276_n 0.00655603f $X=2.24 $Y=2.595 $X2=0 $Y2=0
cc_166 N_A2_c_200_n N_VPWR_c_276_n 0.0101736f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_167 N_A2_M1008_g N_VPWR_c_271_n 0.00846602f $X=2.24 $Y=2.595 $X2=0 $Y2=0
cc_168 N_A2_c_200_n N_VPWR_c_271_n 0.0122683f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_169 N_A2_c_200_n A_359_419# 0.00721535f $X=2.28 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_170 N_A2_c_200_n A_473_419# 0.0110376f $X=2.28 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_171 N_A2_M1004_g N_A_153_57#_c_356_n 0.00776848f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_172 N_A2_M1004_g N_A_153_57#_c_357_n 0.0121208f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_173 N_A2_c_199_n N_A_153_57#_c_357_n 0.00118089f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_174 N_A2_c_200_n N_A_153_57#_c_357_n 0.0194826f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_175 N_A2_M1004_g N_A_153_57#_c_358_n 8.96792e-19 $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_176 N_A2_M1004_g N_A_153_57#_c_359_n 0.00621151f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_177 N_A2_c_200_n N_A_153_57#_c_359_n 0.00632471f $X=2.28 $Y=1.43 $X2=0 $Y2=0
cc_178 N_A2_M1004_g N_VGND_c_411_n 0.00541719f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_179 N_A2_M1004_g N_VGND_c_414_n 0.00502664f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_180 N_A2_M1004_g N_VGND_c_417_n 0.00968694f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_181 N_A1_M1006_g N_VPWR_c_275_n 0.0264908f $X=2.81 $Y=2.595 $X2=0 $Y2=0
cc_182 A1 N_VPWR_c_275_n 0.0278324f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A1_c_244_n N_VPWR_c_275_n 0.00547205f $X=2.975 $Y=1.39 $X2=0 $Y2=0
cc_184 N_A1_M1006_g N_VPWR_c_276_n 0.008763f $X=2.81 $Y=2.595 $X2=0 $Y2=0
cc_185 N_A1_M1006_g N_VPWR_c_271_n 0.0146671f $X=2.81 $Y=2.595 $X2=0 $Y2=0
cc_186 N_A1_M1005_g N_A_153_57#_c_356_n 4.45285e-19 $X=2.78 $Y=0.495 $X2=0 $Y2=0
cc_187 N_A1_M1005_g N_A_153_57#_c_357_n 0.0193012f $X=2.78 $Y=0.495 $X2=0 $Y2=0
cc_188 A1 N_A_153_57#_c_357_n 0.0294073f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A1_c_244_n N_A_153_57#_c_357_n 0.00845987f $X=2.975 $Y=1.39 $X2=0 $Y2=0
cc_190 N_A1_M1005_g N_A_153_57#_c_358_n 0.0128767f $X=2.78 $Y=0.495 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_A_153_57#_c_359_n 4.48261e-19 $X=2.78 $Y=0.495 $X2=0 $Y2=0
cc_192 N_A1_M1005_g N_VGND_c_411_n 0.00541719f $X=2.78 $Y=0.495 $X2=0 $Y2=0
cc_193 N_A1_M1005_g N_VGND_c_416_n 0.00502664f $X=2.78 $Y=0.495 $X2=0 $Y2=0
cc_194 N_A1_M1005_g N_VGND_c_417_n 0.0103741f $X=2.78 $Y=0.495 $X2=0 $Y2=0
cc_195 N_VPWR_c_271_n N_Y_M1002_d 0.00223819f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_M1002_s N_Y_c_313_n 0.00200568f $X=0.23 $Y=2.095 $X2=0 $Y2=0
cc_197 N_VPWR_c_273_n N_Y_c_313_n 0.0151566f $X=0.375 $Y=2.49 $X2=0 $Y2=0
cc_198 N_VPWR_M1002_s N_Y_c_314_n 7.75775e-19 $X=0.23 $Y=2.095 $X2=0 $Y2=0
cc_199 N_VPWR_c_273_n N_Y_c_314_n 0.0064592f $X=0.375 $Y=2.49 $X2=0 $Y2=0
cc_200 N_VPWR_c_273_n N_Y_c_322_n 0.0487591f $X=0.375 $Y=2.49 $X2=0 $Y2=0
cc_201 N_VPWR_c_276_n N_Y_c_322_n 0.0177952f $X=2.91 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_271_n N_Y_c_322_n 0.0123247f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_271_n A_259_419# 0.0107073f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_204 N_VPWR_c_271_n A_359_419# 0.00905433f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_205 N_VPWR_c_271_n A_473_419# 0.0110428f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_206 N_Y_c_310_n N_A_153_57#_c_353_n 0.00175979f $X=0.2 $Y=1.975 $X2=0 $Y2=0
cc_207 N_Y_c_311_n N_A_153_57#_c_353_n 0.0180757f $X=0.395 $Y=0.495 $X2=0 $Y2=0
cc_208 N_Y_c_310_n N_A_153_57#_c_355_n 0.00645337f $X=0.2 $Y=1.975 $X2=0 $Y2=0
cc_209 N_Y_c_311_n N_VGND_c_412_n 0.0293385f $X=0.395 $Y=0.495 $X2=0 $Y2=0
cc_210 N_Y_c_311_n N_VGND_c_417_n 0.0170318f $X=0.395 $Y=0.495 $X2=0 $Y2=0
cc_211 N_A_153_57#_c_353_n N_VGND_c_410_n 0.0125869f $X=0.905 $Y=0.495 $X2=0
+ $Y2=0
cc_212 N_A_153_57#_c_354_n N_VGND_c_410_n 0.025104f $X=1.81 $Y=0.86 $X2=0 $Y2=0
cc_213 N_A_153_57#_c_356_n N_VGND_c_410_n 0.0203419f $X=1.975 $Y=0.495 $X2=0
+ $Y2=0
cc_214 N_A_153_57#_c_356_n N_VGND_c_411_n 0.016171f $X=1.975 $Y=0.495 $X2=0
+ $Y2=0
cc_215 N_A_153_57#_c_357_n N_VGND_c_411_n 0.0259275f $X=2.83 $Y=0.96 $X2=0 $Y2=0
cc_216 N_A_153_57#_c_358_n N_VGND_c_411_n 0.016171f $X=2.995 $Y=0.495 $X2=0
+ $Y2=0
cc_217 N_A_153_57#_c_353_n N_VGND_c_412_n 0.021949f $X=0.905 $Y=0.495 $X2=0
+ $Y2=0
cc_218 N_A_153_57#_c_356_n N_VGND_c_414_n 0.021949f $X=1.975 $Y=0.495 $X2=0
+ $Y2=0
cc_219 N_A_153_57#_c_358_n N_VGND_c_416_n 0.0220321f $X=2.995 $Y=0.495 $X2=0
+ $Y2=0
cc_220 N_A_153_57#_c_353_n N_VGND_c_417_n 0.0124703f $X=0.905 $Y=0.495 $X2=0
+ $Y2=0
cc_221 N_A_153_57#_c_354_n N_VGND_c_417_n 0.0144229f $X=1.81 $Y=0.86 $X2=0 $Y2=0
cc_222 N_A_153_57#_c_356_n N_VGND_c_417_n 0.0124703f $X=1.975 $Y=0.495 $X2=0
+ $Y2=0
cc_223 N_A_153_57#_c_358_n N_VGND_c_417_n 0.0125808f $X=2.995 $Y=0.495 $X2=0
+ $Y2=0
