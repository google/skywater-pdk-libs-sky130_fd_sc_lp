* File: sky130_fd_sc_lp__iso0p_lp2.spice
* Created: Wed Sep  2 09:57:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__iso0p_lp2.pex.spice"
.subckt sky130_fd_sc_lp__iso0p_lp2  VNB VPB SLEEP A KAPWR X VGND VPWR
* 
* VGND	VGND
* X	X
* KAPWR	KAPWR
* A	A
* SLEEP	SLEEP
* VPB	VPB
* VNB	VNB
MM1008 A_112_93# N_SLEEP_M1008_g N_A_27_93#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_SLEEP_M1003_g A_112_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1323 AS=0.0441 PD=1.05 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 A_340_93# N_A_27_93#_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1323 PD=0.63 PS=1.05 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_342_417#_M1000_d N_A_M1000_g A_340_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_602_93# N_A_342_417#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_342_417#_M1002_g A_602_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_KAPWR_M1007_d N_SLEEP_M1007_g N_A_27_93#_M1007_s VPB PHIGHVT L=0.25 W=1
+ AD=0.4 AS=0.275 PD=1.8 PS=2.55 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1009 N_A_342_417#_M1009_d N_A_27_93#_M1009_g N_KAPWR_M1007_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.15 AS=0.4 PD=1.3 PS=1.8 NRD=3.9203 NRS=0 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1005 N_KAPWR_M1005_d N_A_M1005_g N_A_342_417#_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.43 AS=0.15 PD=1.86 PS=1.3 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_X_M1006_d N_A_342_417#_M1006_g N_KAPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.43 PD=2.53 PS=1.86 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.86097 P=12.16
*
.include "sky130_fd_sc_lp__iso0p_lp2.pxi.spice"
*
.ends
*
*
