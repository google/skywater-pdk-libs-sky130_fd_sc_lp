* NGSPICE file created from sky130_fd_sc_lp__nand2_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand2_lp A B VGND VNB VPB VPWR Y
M1000 a_121_57# B VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_207_367# A Y VPB phighvt w=420000u l=150000u
+  ad=2.6835e+11p pd=2.89e+06u as=1.176e+11p ps=1.4e+06u
M1002 VPWR B a_39_367# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.6835e+11p ps=2.89e+06u
M1003 Y B a_39_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A a_121_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1005 a_207_367# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

