* File: sky130_fd_sc_lp__and2_lp2.pex.spice
* Created: Fri Aug 28 10:04:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2_LP2%A_99_21# 1 2 7 9 12 16 19 21 22 23 24 26 27
+ 30 36 40
c69 21 0 1.07716e-19 $X=0.68 $Y=1.485
c70 12 0 3.08033e-20 $X=0.71 $Y=2.545
r71 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7 $Y=0.98
+ $X2=0.7 $Y2=0.98
r72 34 36 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.965 $Y=0.815
+ $X2=1.965 $Y2=0.47
r73 30 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.505 $Y=2.19
+ $X2=1.505 $Y2=2.9
r74 28 30 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.505 $Y=1.845
+ $X2=1.505 $Y2=2.19
r75 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.34 $Y=1.76
+ $X2=1.505 $Y2=1.845
r76 26 27 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.34 $Y=1.76
+ $X2=0.865 $Y2=1.76
r77 25 39 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0.9 $X2=0.7
+ $Y2=0.9
r78 24 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.8 $Y=0.9
+ $X2=1.965 $Y2=0.815
r79 24 25 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.8 $Y=0.9 $X2=0.865
+ $Y2=0.9
r80 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.7 $Y=1.675
+ $X2=0.865 $Y2=1.76
r81 22 39 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.985 $X2=0.7
+ $Y2=0.9
r82 22 23 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=0.7 $Y=0.985 $X2=0.7
+ $Y2=1.675
r83 20 40 49.9064 $w=3.7e-07 $l=3.2e-07 $layer=POLY_cond $X=0.68 $Y=1.3 $X2=0.68
+ $Y2=0.98
r84 20 21 32.9177 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=0.68 $Y=1.3
+ $X2=0.68 $Y2=1.485
r85 19 40 8.57765 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=0.68 $Y=0.925
+ $X2=0.68 $Y2=0.98
r86 12 21 263.361 $w=2.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.71 $Y=2.545
+ $X2=0.71 $Y2=1.485
r87 7 19 25.6283 $w=3.7e-07 $l=1.5e-07 $layer=POLY_cond $X=0.75 $Y=0.775
+ $X2=0.75 $Y2=0.925
r88 7 16 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.93 $Y=0.775 $X2=0.93
+ $Y2=0.445
r89 7 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.57 $Y=0.775 $X2=0.57
+ $Y2=0.445
r90 2 32 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.045 $X2=1.505 $Y2=2.9
r91 2 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.045 $X2=1.505 $Y2=2.19
r92 1 36 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.965 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP2%B 3 7 9 12
c38 9 0 3.08033e-20 $X=1.2 $Y=1.295
r39 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.27 $Y=1.33
+ $X2=1.27 $Y2=1.495
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.27 $Y=1.33
+ $X2=1.27 $Y2=1.165
r41 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.33 $X2=1.27 $Y2=1.33
r42 7 14 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.36 $Y=0.445
+ $X2=1.36 $Y2=1.165
r43 3 15 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.24 $Y=2.545
+ $X2=1.24 $Y2=1.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP2%A 3 7 9 10 14
r29 14 17 67.1496 $w=5.05e-07 $l=5.05e-07 $layer=POLY_cond $X=1.927 $Y=1.33
+ $X2=1.927 $Y2=1.835
r30 14 16 46.6818 $w=5.05e-07 $l=1.65e-07 $layer=POLY_cond $X=1.927 $Y=1.33
+ $X2=1.927 $Y2=1.165
r31 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.015
+ $Y=1.33 $X2=2.015 $Y2=1.33
r32 10 15 9.08396 $w=4.23e-07 $l=3.35e-07 $layer=LI1_cond $X=2.062 $Y=1.665
+ $X2=2.062 $Y2=1.33
r33 9 15 0.949071 $w=4.23e-07 $l=3.5e-08 $layer=LI1_cond $X=2.062 $Y=1.295
+ $X2=2.062 $Y2=1.33
r34 7 17 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.8 $Y=2.545 $X2=1.8
+ $Y2=1.835
r35 3 16 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.75 $Y=0.445
+ $X2=1.75 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP2%X 1 2 7 8 9 10 11 12 13 45 48
r23 48 49 3.57067 $w=4.83e-07 $l=1e-08 $layer=LI1_cond $X=0.367 $Y=2.035
+ $X2=0.367 $Y2=2.025
r24 33 52 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=0.367 $Y=2.267
+ $X2=0.367 $Y2=2.19
r25 13 39 3.08268 $w=4.83e-07 $l=1.25e-07 $layer=LI1_cond $X=0.367 $Y=2.775
+ $X2=0.367 $Y2=2.9
r26 12 13 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.367 $Y=2.405
+ $X2=0.367 $Y2=2.775
r27 12 33 3.40327 $w=4.83e-07 $l=1.38e-07 $layer=LI1_cond $X=0.367 $Y=2.405
+ $X2=0.367 $Y2=2.267
r28 11 52 2.91005 $w=4.83e-07 $l=1.18e-07 $layer=LI1_cond $X=0.367 $Y=2.072
+ $X2=0.367 $Y2=2.19
r29 11 48 0.912472 $w=4.83e-07 $l=3.7e-08 $layer=LI1_cond $X=0.367 $Y=2.072
+ $X2=0.367 $Y2=2.035
r30 11 49 1.90404 $w=2.28e-07 $l=3.8e-08 $layer=LI1_cond $X=0.24 $Y=1.987
+ $X2=0.24 $Y2=2.025
r31 10 11 16.1342 $w=2.28e-07 $l=3.22e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.987
r32 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r33 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925 $X2=0.24
+ $Y2=1.295
r34 7 45 3.58192 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=0.45
+ $X2=0.355 $Y2=0.45
r35 7 23 3.51871 $w=2.3e-07 $l=1.85e-07 $layer=LI1_cond $X=0.24 $Y=0.45 $X2=0.24
+ $Y2=0.635
r36 7 8 14.4306 $w=2.28e-07 $l=2.88e-07 $layer=LI1_cond $X=0.24 $Y=0.637
+ $X2=0.24 $Y2=0.925
r37 7 23 0.100212 $w=2.28e-07 $l=2e-09 $layer=LI1_cond $X=0.24 $Y=0.637 $X2=0.24
+ $Y2=0.635
r38 2 52 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=2.045 $X2=0.445 $Y2=2.19
r39 2 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=2.045 $X2=0.445 $Y2=2.9
r40 1 45 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.21
+ $Y=0.235 $X2=0.355 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP2%VPWR 1 2 9 13 15 20 21 22 28 34
c30 9 0 1.07716e-19 $X=0.975 $Y=2.19
r31 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 28 33 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.9 $Y=3.33 $X2=2.15
+ $Y2=3.33
r35 28 30 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.9 $Y=3.33 $X2=1.68
+ $Y2=3.33
r36 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 22 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 20 25 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.81 $Y=3.33 $X2=0.72
+ $Y2=3.33
r40 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=3.33
+ $X2=0.975 $Y2=3.33
r41 19 30 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.14 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=3.33
+ $X2=0.975 $Y2=3.33
r43 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.065 $Y=2.19
+ $X2=2.065 $Y2=2.9
r44 13 33 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=3.245
+ $X2=2.15 $Y2=3.33
r45 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.065 $Y=3.245
+ $X2=2.065 $Y2=2.9
r46 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.975 $Y=2.19
+ $X2=0.975 $Y2=2.9
r47 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=3.245
+ $X2=0.975 $Y2=3.33
r48 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.975 $Y=3.245
+ $X2=0.975 $Y2=2.9
r49 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=2.045 $X2=2.065 $Y2=2.9
r50 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=2.045 $X2=2.065 $Y2=2.19
r51 1 12 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.835
+ $Y=2.045 $X2=0.975 $Y2=2.9
r52 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.835
+ $Y=2.045 $X2=0.975 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP2%VGND 1 6 8 10 17 18 21
r29 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r30 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=1.145
+ $Y2=0
r31 15 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=2.16
+ $Y2=0
r32 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.145
+ $Y2=0
r34 10 12 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.72
+ $Y2=0
r35 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r36 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r37 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0
r39 4 6 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0.425
r40 1 6 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.145 $Y2=0.425
.ends

