* File: sky130_fd_sc_lp__xnor2_m.spice
* Created: Wed Sep  2 10:40:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor2_m.pex.spice"
.subckt sky130_fd_sc_lp__xnor2_m  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_139_90# N_B_M1002_g N_A_56_90#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g A_139_90# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_297_90#_M1003_d N_A_M1003_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g N_A_297_90#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0588 PD=1.53 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1006 N_A_297_90#_M1006_d N_A_56_90#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_56_90#_M1000_d N_B_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_56_90#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1008 A_311_422# N_A_M1008_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g A_311_422# VPB PHIGHVT L=0.15 W=0.42 AD=0.1575
+ AS=0.0441 PD=1.17 PS=0.63 NRD=157.127 NRS=23.443 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_56_90#_M1004_g N_Y_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.126 AS=0.1575 PD=1.44 PS=1.17 NRD=16.4101 NRS=63.3158 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_59 VPB 0 1.45309e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__xnor2_m.pxi.spice"
*
.ends
*
*
