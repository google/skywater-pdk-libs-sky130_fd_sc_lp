* File: sky130_fd_sc_lp__nand2b_2.pex.spice
* Created: Wed Sep  2 10:03:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2B_2%A_N 1 3 4 6 8
c29 1 0 1.30779e-19 $X=0.475 $Y=1.185
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.35 $X2=0.525 $Y2=1.35
r31 8 12 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.72 $Y=1.35
+ $X2=0.525 $Y2=1.35
r32 4 11 38.6287 $w=3.34e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.625 $Y=1.515
+ $X2=0.53 $Y2=1.35
r33 4 6 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.625 $Y=1.515
+ $X2=0.625 $Y2=2.045
r34 1 11 38.6287 $w=3.34e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.53 $Y2=1.35
r35 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_2%B 3 6 10 13 15 17 21 23 26 28 31 33
c78 26 0 1.15358e-19 $X=1.095 $Y=1.35
r79 26 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.35
+ $X2=1.095 $Y2=1.515
r80 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.35
+ $X2=1.095 $Y2=1.185
r81 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.35 $X2=1.095 $Y2=1.35
r82 23 27 2.18567 $w=2.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.35
r83 23 33 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.16
r84 21 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.53 $Y=1.35
+ $X2=2.53 $Y2=1.515
r85 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.53 $Y=1.35
+ $X2=2.53 $Y2=1.185
r86 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.35 $X2=2.53 $Y2=1.35
r87 17 20 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.53 $Y=1.16
+ $X2=2.53 $Y2=1.35
r88 16 33 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.3 $Y=1.16
+ $X2=1.155 $Y2=1.16
r89 15 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=1.16
+ $X2=2.53 $Y2=1.16
r90 15 16 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=2.365 $Y=1.16
+ $X2=1.3 $Y2=1.16
r91 13 32 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.44 $Y=2.465
+ $X2=2.44 $Y2=1.515
r92 10 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.44 $Y=0.655
+ $X2=2.44 $Y2=1.185
r93 6 29 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.15 $Y=2.465
+ $X2=1.15 $Y2=1.515
r94 3 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.07 $Y=0.655
+ $X2=1.07 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_2%A_27_131# 1 2 9 13 17 21 25 30 32 33 38 47
c74 38 0 1.15358e-19 $X=1.635 $Y=1.51
r75 43 45 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.545 $Y=1.51
+ $X2=1.58 $Y2=1.51
r76 39 47 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.635 $Y=1.51
+ $X2=2.01 $Y2=1.51
r77 39 45 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.635 $Y=1.51
+ $X2=1.58 $Y2=1.51
r78 38 41 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.635 $Y=1.51
+ $X2=1.635 $Y2=1.78
r79 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.51 $X2=1.635 $Y2=1.51
r80 32 35 7.35897 $w=4.13e-07 $l=2.65e-07 $layer=LI1_cond $X=0.297 $Y=1.78
+ $X2=0.297 $Y2=2.045
r81 32 33 6.49176 $w=4.13e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=1.78
+ $X2=0.297 $Y2=1.695
r82 27 30 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.175 $Y=0.85
+ $X2=0.26 $Y2=0.85
r83 26 32 6.00275 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.505 $Y=1.78
+ $X2=0.297 $Y2=1.78
r84 25 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=1.78
+ $X2=1.635 $Y2=1.78
r85 25 26 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.47 $Y=1.78
+ $X2=0.505 $Y2=1.78
r86 23 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.175 $Y=1.015
+ $X2=0.175 $Y2=0.85
r87 23 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.175 $Y=1.015
+ $X2=0.175 $Y2=1.695
r88 19 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.675
+ $X2=2.01 $Y2=1.51
r89 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.01 $Y=1.675
+ $X2=2.01 $Y2=2.465
r90 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.345
+ $X2=2.01 $Y2=1.51
r91 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.01 $Y=1.345
+ $X2=2.01 $Y2=0.655
r92 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.675
+ $X2=1.58 $Y2=1.51
r93 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.58 $Y=1.675
+ $X2=1.58 $Y2=2.465
r94 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.545 $Y=1.345
+ $X2=1.545 $Y2=1.51
r95 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.545 $Y=1.345
+ $X2=1.545 $Y2=0.655
r96 2 35 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.835 $X2=0.41 $Y2=2.045
r97 1 30 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.655 $X2=0.26 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_2%VPWR 1 2 3 14 18 22 26 28 30 37 38 41 44 47
r40 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 38 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 35 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.655 $Y2=3.33
r45 35 37 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.82 $Y=3.33 $X2=3.12
+ $Y2=3.33
r46 34 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.96 $Y=3.33
+ $X2=1.795 $Y2=3.33
r49 31 33 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.96 $Y=3.33 $X2=2.16
+ $Y2=3.33
r50 30 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.655 $Y2=3.33
r51 30 33 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 28 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 28 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 24 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.655 $Y=3.245
+ $X2=2.655 $Y2=3.33
r56 24 26 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.655 $Y=3.245
+ $X2=2.655 $Y2=2.41
r57 20 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=3.245
+ $X2=1.795 $Y2=3.33
r58 20 22 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.795 $Y=3.245
+ $X2=1.795 $Y2=2.485
r59 19 41 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.867 $Y2=3.33
r60 18 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=3.33
+ $X2=1.795 $Y2=3.33
r61 18 19 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.63 $Y=3.33
+ $X2=1.06 $Y2=3.33
r62 14 17 12.7218 $w=3.83e-07 $l=4.25e-07 $layer=LI1_cond $X=0.867 $Y=2.12
+ $X2=0.867 $Y2=2.545
r63 12 41 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.867 $Y=3.245
+ $X2=0.867 $Y2=3.33
r64 12 17 20.9535 $w=3.83e-07 $l=7e-07 $layer=LI1_cond $X=0.867 $Y=3.245
+ $X2=0.867 $Y2=2.545
r65 3 26 300 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=1.835 $X2=2.655 $Y2=2.41
r66 2 22 300 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=2 $X=1.655
+ $Y=1.835 $X2=1.795 $Y2=2.485
r67 1 17 300 $w=1.7e-07 $l=8.19115e-07 $layer=licon1_PDIFF $count=2 $X=0.7
+ $Y=1.835 $X2=0.935 $Y2=2.545
r68 1 14 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.7
+ $Y=1.835 $X2=0.84 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_2%Y 1 2 3 10 12 16 20 23 29 30 31 32 36 41 44
r50 32 36 4.08363 $w=2.9e-07 $l=2e-07 $layer=LI1_cond $X=3.075 $Y=1.975
+ $X2=2.875 $Y2=1.975
r51 31 36 9.33876 $w=2.88e-07 $l=2.35e-07 $layer=LI1_cond $X=2.64 $Y=1.975
+ $X2=2.875 $Y2=1.975
r52 31 44 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=2.64 $Y=1.975
+ $X2=2.32 $Y2=1.975
r53 30 44 5.5393 $w=3.73e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=2.017
+ $X2=2.32 $Y2=2.017
r54 30 41 9.32276 $w=3.73e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=2.017
+ $X2=1.97 $Y2=2.017
r55 27 29 8.52828 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0.78
+ $X2=1.96 $Y2=0.78
r56 23 32 2.96063 $w=4e-07 $l=1.45e-07 $layer=LI1_cond $X=3.075 $Y=1.83
+ $X2=3.075 $Y2=1.975
r57 22 23 26.6502 $w=3.98e-07 $l=9.25e-07 $layer=LI1_cond $X=3.075 $Y=0.905
+ $X2=3.075 $Y2=1.83
r58 18 30 4.72237 $w=1.9e-07 $l=2.18092e-07 $layer=LI1_cond $X=2.225 $Y=2.205
+ $X2=2.16 $Y2=2.017
r59 18 20 14.0096 $w=1.88e-07 $l=2.4e-07 $layer=LI1_cond $X=2.225 $Y=2.205
+ $X2=2.225 $Y2=2.445
r60 16 22 8.17735 $w=1.8e-07 $l=2.40832e-07 $layer=LI1_cond $X=2.875 $Y=0.815
+ $X2=3.075 $Y2=0.905
r61 16 29 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=2.875 $Y=0.815
+ $X2=1.96 $Y2=0.815
r62 15 25 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.46 $Y=2.12
+ $X2=1.345 $Y2=2.12
r63 15 41 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.46 $Y=2.12
+ $X2=1.97 $Y2=2.12
r64 10 25 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.345 $Y=2.205
+ $X2=1.345 $Y2=2.12
r65 10 12 35.3249 $w=2.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.345 $Y=2.205
+ $X2=1.345 $Y2=2.91
r66 3 30 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=1.835 $X2=2.225 $Y2=1.995
r67 3 20 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=2.085
+ $Y=1.835 $X2=2.225 $Y2=2.445
r68 2 25 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=1.835 $X2=1.365 $Y2=2.2
r69 2 12 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=1.835 $X2=1.365 $Y2=2.91
r70 1 27 182 $w=1.7e-07 $l=6.36514e-07 $layer=licon1_NDIFF $count=1 $X=1.62
+ $Y=0.235 $X2=1.795 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_2%VGND 1 2 8 10 13 17 19 24 31 32 35 38
r41 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r44 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 29 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=2.69
+ $Y2=0
r46 29 31 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=3.12
+ $Y2=0
r47 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 25 35 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.737
+ $Y2=0
r50 25 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r51 24 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.69
+ $Y2=0
r52 24 27 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=0 $X2=1.2
+ $Y2=0
r53 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 19 35 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.737
+ $Y2=0
r56 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r57 17 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r58 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 11 38 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=0.085
+ $X2=2.69 $Y2=0
r60 11 13 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.69 $Y=0.085
+ $X2=2.69 $Y2=0.39
r61 8 16 4.5814 $w=4.25e-07 $l=1.57e-07 $layer=LI1_cond $X=0.737 $Y=0.693
+ $X2=0.737 $Y2=0.85
r62 8 10 8.4874 $w=4.23e-07 $l=3.13e-07 $layer=LI1_cond $X=0.737 $Y=0.693
+ $X2=0.737 $Y2=0.38
r63 7 35 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0
r64 7 10 7.99931 $w=4.23e-07 $l=2.95e-07 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0.38
r65 2 13 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.235 $X2=2.655 $Y2=0.39
r66 1 16 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.655 $X2=0.69 $Y2=0.85
r67 1 10 182 $w=1.7e-07 $l=4.20595e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.655 $X2=0.855 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_2%A_229_47# 1 2 7 9 13
c20 9 0 1.30779e-19 $X=1.285 $Y=0.82
r21 11 16 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0.37
+ $X2=1.285 $Y2=0.37
r22 11 13 38.8323 $w=2.28e-07 $l=7.75e-07 $layer=LI1_cond $X=1.45 $Y=0.37
+ $X2=2.225 $Y2=0.37
r23 7 16 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.285 $Y=0.485
+ $X2=1.285 $Y2=0.37
r24 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.285 $Y=0.485
+ $X2=1.285 $Y2=0.82
r25 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.225 $Y2=0.38
r26 1 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.235 $X2=1.285 $Y2=0.38
r27 1 9 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.235 $X2=1.285 $Y2=0.82
.ends

