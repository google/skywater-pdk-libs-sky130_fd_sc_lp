* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_151_367# A3 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=8.883e+11p ps=6.45e+06u
M1001 a_151_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=4.494e+11p pd=4.43e+06u as=3.276e+11p ps=2.46e+06u
M1003 a_151_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1004 Y B1 a_151_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.347e+11p pd=3.21e+06u as=0p ps=0u
M1005 VPWR A2 a_151_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_223_47# A2 a_151_47# VNB nshort w=840000u l=150000u
+  ad=3.36e+11p pd=2.48e+06u as=0p ps=0u
M1007 Y A1 a_223_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
