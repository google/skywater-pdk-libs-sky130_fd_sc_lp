* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__inv_8 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=1.7766e+12p pd=1.542e+07u as=1.4112e+12p ps=1.232e+07u
M1001 VGND A Y VNB nshort w=840000u l=150000u
+  ad=1.1844e+12p pd=1.122e+07u as=9.408e+11p ps=8.96e+06u
M1002 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
