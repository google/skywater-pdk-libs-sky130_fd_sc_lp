* File: sky130_fd_sc_lp__mux4_4.pex.spice
* Created: Fri Aug 28 10:46:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX4_4%A_84_277# 1 2 9 11 12 15 17 19 22 27 28 29 34
r56 31 34 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=0.805
+ $X2=1.94 $Y2=0.805
r57 28 38 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.51 $Y=1.315
+ $X2=1.51 $Y2=1.46
r58 27 30 13.9269 $w=4.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.66 $Y=1.315
+ $X2=1.66 $Y2=1.82
r59 27 29 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.315
+ $X2=1.66 $Y2=1.15
r60 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.51
+ $Y=1.315 $X2=1.51 $Y2=1.315
r61 24 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=0.97
+ $X2=1.81 $Y2=0.805
r62 24 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.81 $Y=0.97
+ $X2=1.81 $Y2=1.15
r63 22 30 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.73 $Y=2.105
+ $X2=1.73 $Y2=1.82
r64 18 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1 $Y=1.46 $X2=0.925
+ $Y2=1.46
r65 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.46
+ $X2=1.51 $Y2=1.46
r66 17 18 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.345 $Y=1.46 $X2=1
+ $Y2=1.46
r67 13 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.925 $Y=1.385
+ $X2=0.925 $Y2=1.46
r68 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.925 $Y=1.385
+ $X2=0.925 $Y2=0.805
r69 11 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.85 $Y=1.46
+ $X2=0.925 $Y2=1.46
r70 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.85 $Y=1.46
+ $X2=0.57 $Y2=1.46
r71 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=1.535
+ $X2=0.57 $Y2=1.46
r72 7 9 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.495 $Y=1.535
+ $X2=0.495 $Y2=2.33
r73 2 22 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=1.98 $X2=1.73 $Y2=2.105
r74 1 34 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.655 $X2=1.94 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%S1 3 5 6 7 9 10 11 15 19 20 21 22 27
r69 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.35
+ $X2=2.16 $Y2=1.185
r70 21 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=2.035
r71 20 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r72 20 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.35 $X2=2.16 $Y2=1.35
r73 19 29 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.175 $Y=0.865
+ $X2=2.175 $Y2=1.185
r74 16 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.175 $Y=0.255
+ $X2=2.175 $Y2=0.865
r75 13 15 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.16 $Y=2.76
+ $X2=2.16 $Y2=1.995
r76 12 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.515
+ $X2=2.16 $Y2=1.35
r77 12 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.16 $Y=1.515
+ $X2=2.16 $Y2=1.995
r78 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.085 $Y=2.835
+ $X2=2.16 $Y2=2.76
r79 10 11 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=2.085 $Y=2.835
+ $X2=1 $Y2=2.835
r80 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=2.76
+ $X2=1 $Y2=2.835
r81 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.925 $Y=2.76
+ $X2=0.925 $Y2=2.33
r82 5 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.1 $Y=0.18
+ $X2=2.175 $Y2=0.255
r83 5 6 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=2.1 $Y=0.18 $X2=0.57
+ $Y2=0.18
r84 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.57 $Y2=0.18
r85 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.495 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A_114_119# 1 2 9 11 13 16 18 20 23 25 27 30
+ 32 34 37 41 42 44 45 46 48 49 54 65
c135 65 0 1.14729e-19 $X=3.995 $Y=1.35
r136 64 65 43.1182 $w=3.13e-07 $l=2.8e-07 $layer=POLY_cond $X=3.715 $Y=1.35
+ $X2=3.995 $Y2=1.35
r137 63 64 23.099 $w=3.13e-07 $l=1.5e-07 $layer=POLY_cond $X=3.565 $Y=1.35
+ $X2=3.715 $Y2=1.35
r138 60 61 23.099 $w=3.13e-07 $l=1.5e-07 $layer=POLY_cond $X=3.135 $Y=1.35
+ $X2=3.285 $Y2=1.35
r139 59 60 43.1182 $w=3.13e-07 $l=2.8e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=3.135 $Y2=1.35
r140 55 63 13.8594 $w=3.13e-07 $l=9e-08 $layer=POLY_cond $X=3.475 $Y=1.35
+ $X2=3.565 $Y2=1.35
r141 55 61 29.2588 $w=3.13e-07 $l=1.9e-07 $layer=POLY_cond $X=3.475 $Y=1.35
+ $X2=3.285 $Y2=1.35
r142 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.475
+ $Y=1.35 $X2=3.475 $Y2=1.35
r143 52 59 9.23962 $w=3.13e-07 $l=6e-08 $layer=POLY_cond $X=2.795 $Y=1.35
+ $X2=2.855 $Y2=1.35
r144 52 57 13.8594 $w=3.13e-07 $l=9e-08 $layer=POLY_cond $X=2.795 $Y=1.35
+ $X2=2.705 $Y2=1.35
r145 51 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.795 $Y=1.35
+ $X2=3.475 $Y2=1.35
r146 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.35 $X2=2.795 $Y2=1.35
r147 49 51 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.785 $Y=1.35
+ $X2=2.795 $Y2=1.35
r148 48 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.7 $Y=1.265
+ $X2=2.785 $Y2=1.35
r149 47 48 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.7 $Y=1.005
+ $X2=2.7 $Y2=1.265
r150 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.615 $Y=0.92
+ $X2=2.7 $Y2=1.005
r151 45 46 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.615 $Y=0.92
+ $X2=2.375 $Y2=0.92
r152 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.29 $Y=0.835
+ $X2=2.375 $Y2=0.92
r153 43 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.29 $Y=0.46
+ $X2=2.29 $Y2=0.835
r154 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=0.375
+ $X2=2.29 $Y2=0.46
r155 41 42 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.205 $Y=0.375
+ $X2=0.795 $Y2=0.375
r156 37 39 82.5981 $w=1.88e-07 $l=1.415e-06 $layer=LI1_cond $X=0.7 $Y=0.74
+ $X2=0.7 $Y2=2.155
r157 35 42 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.7 $Y=0.46
+ $X2=0.795 $Y2=0.375
r158 35 37 16.3445 $w=1.88e-07 $l=2.8e-07 $layer=LI1_cond $X=0.7 $Y=0.46 $X2=0.7
+ $Y2=0.74
r159 32 65 23.099 $w=3.13e-07 $l=2.2798e-07 $layer=POLY_cond $X=4.145 $Y=1.185
+ $X2=3.995 $Y2=1.35
r160 32 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.145 $Y=1.185
+ $X2=4.145 $Y2=0.655
r161 28 65 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.515
+ $X2=3.995 $Y2=1.35
r162 28 30 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.995 $Y=1.515
+ $X2=3.995 $Y2=2.305
r163 25 64 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.715 $Y=1.185
+ $X2=3.715 $Y2=1.35
r164 25 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.715 $Y=1.185
+ $X2=3.715 $Y2=0.655
r165 21 63 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.515
+ $X2=3.565 $Y2=1.35
r166 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.565 $Y=1.515
+ $X2=3.565 $Y2=2.305
r167 18 61 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.185
+ $X2=3.285 $Y2=1.35
r168 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.285 $Y=1.185
+ $X2=3.285 $Y2=0.655
r169 14 60 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.135 $Y=1.515
+ $X2=3.135 $Y2=1.35
r170 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.135 $Y=1.515
+ $X2=3.135 $Y2=2.305
r171 11 59 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.185
+ $X2=2.855 $Y2=1.35
r172 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.855 $Y=1.185
+ $X2=2.855 $Y2=0.655
r173 7 57 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.515
+ $X2=2.705 $Y2=1.35
r174 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.705 $Y=1.515
+ $X2=2.705 $Y2=2.305
r175 2 39 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.01 $X2=0.71 $Y2=2.155
r176 1 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.595 $X2=0.71 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A1 3 7 9 10 16
c45 16 0 2.38611e-19 $X=4.685 $Y=1.36
c46 7 0 1.6982e-19 $X=4.92 $Y=2.475
r47 14 16 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=4.595 $Y=1.36
+ $X2=4.685 $Y2=1.36
r48 9 10 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=4.577 $Y=1.295
+ $X2=4.577 $Y2=1.665
r49 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.595
+ $Y=1.35 $X2=4.595 $Y2=1.35
r50 5 16 42.5827 $w=2.66e-07 $l=3.10403e-07 $layer=POLY_cond $X=4.92 $Y=1.535
+ $X2=4.685 $Y2=1.36
r51 5 7 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.92 $Y=1.535 $X2=4.92
+ $Y2=2.475
r52 1 16 16.1576 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.685 $Y=1.185
+ $X2=4.685 $Y2=1.36
r53 1 3 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.685 $Y=1.185
+ $X2=4.685 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A_1041_333# 1 2 9 13 17 21 25 28 29 30 33 34
+ 36 39 40 41 44 46 48 55 56 63
c145 63 0 1.93349e-19 $X=5.475 $Y=1.65
c146 55 0 1.09216e-19 $X=7.57 $Y=1.29
c147 41 0 8.13193e-20 $X=8.615 $Y=2.06
c148 33 0 1.98209e-19 $X=7.57 $Y=1.63
r149 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=1.29 $X2=7.57 $Y2=1.29
r150 53 63 37.5471 $w=2.76e-07 $l=2.15e-07 $layer=POLY_cond $X=5.69 $Y=1.65
+ $X2=5.475 $Y2=1.65
r151 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.69
+ $Y=1.65 $X2=5.69 $Y2=1.65
r152 46 48 38.5894 $w=3.28e-07 $l=1.105e-06 $layer=LI1_cond $X=9.33 $Y=1.975
+ $X2=9.33 $Y2=0.87
r153 42 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.025 $Y=2.06
+ $X2=9.33 $Y2=2.06
r154 42 44 5.01732 $w=2.08e-07 $l=9.5e-08 $layer=LI1_cond $X=9.025 $Y=2.145
+ $X2=9.025 $Y2=2.24
r155 40 42 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.92 $Y=2.06
+ $X2=9.025 $Y2=2.06
r156 40 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.92 $Y=2.06
+ $X2=8.615 $Y2=2.06
r157 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.53 $Y=1.975
+ $X2=8.615 $Y2=2.06
r158 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.53 $Y=1.295
+ $X2=8.53 $Y2=1.975
r159 37 55 5.16603 $w=1.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.655 $Y=1.21
+ $X2=7.57 $Y2=1.262
r160 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.445 $Y=1.21
+ $X2=8.53 $Y2=1.295
r161 36 37 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.445 $Y=1.21
+ $X2=7.655 $Y2=1.21
r162 34 56 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.57 $Y=1.63
+ $X2=7.57 $Y2=1.29
r163 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=1.63 $X2=7.57 $Y2=1.63
r164 31 55 1.34256 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=7.57 $Y=1.4
+ $X2=7.57 $Y2=1.262
r165 31 33 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.57 $Y=1.4
+ $X2=7.57 $Y2=1.63
r166 30 52 12.6925 $w=3.22e-07 $l=4.3119e-07 $layer=LI1_cond $X=6.045 $Y=1.315
+ $X2=5.825 $Y2=1.65
r167 29 55 5.16603 $w=1.7e-07 $l=1.08305e-07 $layer=LI1_cond $X=7.485 $Y=1.315
+ $X2=7.57 $Y2=1.262
r168 29 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.485 $Y=1.315
+ $X2=6.045 $Y2=1.315
r169 28 56 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.57 $Y=1.125
+ $X2=7.57 $Y2=1.29
r170 25 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.57 $Y=1.645
+ $X2=7.57 $Y2=1.63
r171 22 25 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.3 $Y=1.72
+ $X2=7.57 $Y2=1.72
r172 21 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.55 $Y=0.805
+ $X2=7.55 $Y2=1.125
r173 15 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.3 $Y=1.795
+ $X2=7.3 $Y2=1.72
r174 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.3 $Y=1.795
+ $X2=7.3 $Y2=2.415
r175 11 63 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.485
+ $X2=5.475 $Y2=1.65
r176 11 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.475 $Y=1.485
+ $X2=5.475 $Y2=0.805
r177 7 63 34.0543 $w=2.76e-07 $l=2.64953e-07 $layer=POLY_cond $X=5.28 $Y=1.815
+ $X2=5.475 $Y2=1.65
r178 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.28 $Y=1.815
+ $X2=5.28 $Y2=2.475
r179 2 44 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.885
+ $Y=2.095 $X2=9.025 $Y2=2.24
r180 1 48 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=9.17
+ $Y=0.595 $X2=9.33 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A0 1 3 4 5 10 12 15 17
c42 17 0 7.35671e-20 $X=6.31 $Y=1.58
c43 12 0 1.93349e-19 $X=6.48 $Y=1.665
r44 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.31 $Y=1.745
+ $X2=6.31 $Y2=1.91
r45 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.31 $Y=1.745
+ $X2=6.31 $Y2=1.58
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=1.745 $X2=6.31 $Y2=1.745
r47 12 16 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.48 $Y=1.745
+ $X2=6.31 $Y2=1.745
r48 10 18 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.22 $Y=2.415
+ $X2=6.22 $Y2=1.91
r49 6 17 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=6.22 $Y=1.275
+ $X2=6.22 $Y2=1.58
r50 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.145 $Y=1.2
+ $X2=6.22 $Y2=1.275
r51 4 5 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.145 $Y=1.2 $X2=5.91
+ $Y2=1.2
r52 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.835 $Y=1.125
+ $X2=5.91 $Y2=1.2
r53 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.835 $Y=1.125
+ $X2=5.835 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A3 3 7 9 12
c37 12 0 1.98209e-19 $X=6.85 $Y=1.745
r38 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.85 $Y=1.745
+ $X2=6.85 $Y2=1.91
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.85 $Y=1.745
+ $X2=6.85 $Y2=1.58
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.745 $X2=6.85 $Y2=1.745
r41 9 13 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=6.96 $Y=1.745
+ $X2=6.85 $Y2=1.745
r42 7 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.94 $Y=2.415
+ $X2=6.94 $Y2=1.91
r43 3 14 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=6.76 $Y=0.805
+ $X2=6.76 $Y2=1.58
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A2 3 7 9 10 11 12 19 20
r45 19 21 31.6066 $w=3.05e-07 $l=2e-07 $layer=POLY_cond $X=8.18 $Y=1.65 $X2=8.38
+ $Y2=1.65
r46 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.18
+ $Y=1.65 $X2=8.18 $Y2=1.65
r47 17 19 25.2852 $w=3.05e-07 $l=1.6e-07 $layer=POLY_cond $X=8.02 $Y=1.65
+ $X2=8.18 $Y2=1.65
r48 11 12 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.05 $Y=2.405
+ $X2=8.05 $Y2=2.775
r49 10 11 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.05 $Y=2.035
+ $X2=8.05 $Y2=2.405
r50 9 10 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.05 $Y=1.665
+ $X2=8.05 $Y2=2.035
r51 9 20 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.05 $Y=1.665
+ $X2=8.05 $Y2=1.65
r52 5 21 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.38 $Y=1.815
+ $X2=8.38 $Y2=1.65
r53 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.38 $Y=1.815 $X2=8.38
+ $Y2=2.415
r54 1 17 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.02 $Y=1.485
+ $X2=8.02 $Y2=1.65
r55 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.02 $Y=1.485 $X2=8.02
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%S0 3 5 6 9 11 12 15 17 21 23 26 30 34 35 36
+ 37 38 39 40 41 47
c110 21 0 8.13193e-20 $X=7.87 $Y=2.475
c111 15 0 1.09216e-19 $X=7.12 $Y=0.805
r112 47 49 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=8.952 $Y=1.29
+ $X2=8.952 $Y2=1.125
r113 40 41 21.89 $w=1.88e-07 $l=3.75e-07 $layer=LI1_cond $X=8.89 $Y=1.29
+ $X2=8.89 $Y2=1.665
r114 40 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.9
+ $Y=1.29 $X2=8.9 $Y2=1.29
r115 39 40 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=8.89 $Y=0.925
+ $X2=8.89 $Y2=1.29
r116 38 39 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=8.89 $Y=0.555
+ $X2=8.89 $Y2=0.925
r117 34 49 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.095 $Y=0.805
+ $X2=9.095 $Y2=1.125
r118 31 34 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=9.095 $Y=0.255
+ $X2=9.095 $Y2=0.805
r119 30 37 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.81 $Y=2.415
+ $X2=8.81 $Y2=1.795
r120 28 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.81 $Y=3.075
+ $X2=8.81 $Y2=2.415
r121 26 37 53.1843 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=8.952 $Y=1.578
+ $X2=8.952 $Y2=1.795
r122 25 47 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=8.952 $Y=1.342
+ $X2=8.952 $Y2=1.29
r123 25 26 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=8.952 $Y=1.342
+ $X2=8.952 $Y2=1.578
r124 24 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.945 $Y=3.15
+ $X2=7.87 $Y2=3.15
r125 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.735 $Y=3.15
+ $X2=8.81 $Y2=3.075
r126 23 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.735 $Y=3.15
+ $X2=7.945 $Y2=3.15
r127 19 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.87 $Y=3.075
+ $X2=7.87 $Y2=3.15
r128 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.87 $Y=3.075 $X2=7.87
+ $Y2=2.475
r129 18 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.195 $Y=0.18
+ $X2=7.12 $Y2=0.18
r130 17 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.02 $Y=0.18
+ $X2=9.095 $Y2=0.255
r131 17 18 935.798 $w=1.5e-07 $l=1.825e-06 $layer=POLY_cond $X=9.02 $Y=0.18
+ $X2=7.195 $Y2=0.18
r132 13 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.12 $Y=0.255
+ $X2=7.12 $Y2=0.18
r133 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.12 $Y=0.255
+ $X2=7.12 $Y2=0.805
r134 11 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.795 $Y=3.15
+ $X2=7.87 $Y2=3.15
r135 11 12 1030.66 $w=1.5e-07 $l=2.01e-06 $layer=POLY_cond $X=7.795 $Y=3.15
+ $X2=5.785 $Y2=3.15
r136 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.71 $Y=3.075
+ $X2=5.785 $Y2=3.15
r137 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.71 $Y=3.075 $X2=5.71
+ $Y2=2.475
r138 5 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.045 $Y=0.18
+ $X2=7.12 $Y2=0.18
r139 5 6 987.074 $w=1.5e-07 $l=1.925e-06 $layer=POLY_cond $X=7.045 $Y=0.18
+ $X2=5.12 $Y2=0.18
r140 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.045 $Y=0.255
+ $X2=5.12 $Y2=0.18
r141 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.045 $Y=0.255
+ $X2=5.045 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A_27_119# 1 2 3 4 14 15 16 17 18 19 24 29 30
+ 31 34 37 38
c165 18 0 7.35671e-20 $X=5.695 $Y=0.965
c166 17 0 4.44719e-20 $X=6.475 $Y=0.965
c167 16 0 3.17558e-19 $X=5.425 $Y=2.175
r168 43 45 74.7316 $w=2.08e-07 $l=1.415e-06 $layer=LI1_cond $X=0.26 $Y=0.74
+ $X2=0.26 $Y2=2.155
r169 38 50 7.22718 $w=2.93e-07 $l=1.85e-07 $layer=LI1_cond $X=7.377 $Y=0.555
+ $X2=7.377 $Y2=0.74
r170 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0.555
+ $X2=7.44 $Y2=0.555
r171 34 43 9.77056 $w=2.08e-07 $l=1.85e-07 $layer=LI1_cond $X=0.26 $Y=0.555
+ $X2=0.26 $Y2=0.74
r172 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0.555
+ $X2=0.24 $Y2=0.555
r173 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=0.555
+ $X2=0.24 $Y2=0.555
r174 30 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=0.555
+ $X2=7.44 $Y2=0.555
r175 30 31 8.55196 $w=1.4e-07 $l=6.91e-06 $layer=MET1_cond $X=7.295 $Y=0.555
+ $X2=0.385 $Y2=0.555
r176 24 26 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.56 $Y=0.82
+ $X2=6.56 $Y2=0.965
r177 20 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=0.82
+ $X2=6.56 $Y2=0.82
r178 19 50 3.12527 $w=2.93e-07 $l=8e-08 $layer=LI1_cond $X=7.377 $Y=0.82
+ $X2=7.377 $Y2=0.74
r179 19 20 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=7.23 $Y=0.82
+ $X2=6.645 $Y2=0.82
r180 18 23 17.785 $w=2.68e-07 $l=4.31712e-07 $layer=LI1_cond $X=5.695 $Y=0.965
+ $X2=5.34 $Y2=1.135
r181 17 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=0.965
+ $X2=6.56 $Y2=0.965
r182 17 18 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.475 $Y=0.965
+ $X2=5.695 $Y2=0.965
r183 15 29 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.41 $Y=2.175
+ $X2=7.515 $Y2=2.175
r184 15 16 129.503 $w=1.68e-07 $l=1.985e-06 $layer=LI1_cond $X=7.41 $Y=2.175
+ $X2=5.425 $Y2=2.175
r185 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.34 $Y=2.09
+ $X2=5.425 $Y2=2.175
r186 13 23 3.40055 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.34 $Y=1.305
+ $X2=5.34 $Y2=1.135
r187 13 14 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=5.34 $Y=1.305
+ $X2=5.34 $Y2=2.09
r188 4 29 300 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=2 $X=7.375
+ $Y=2.095 $X2=7.515 $Y2=2.255
r189 3 45 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.01 $X2=0.26 $Y2=2.155
r190 2 50 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.595 $X2=7.335 $Y2=0.74
r191 1 43 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.595 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%A_200_119# 1 2 3 4 13 15 19 22 23 24 26 28 29
+ 31 38 40
c102 40 0 8.77531e-20 $X=4.99 $Y=2.08
c103 38 0 1.71397e-19 $X=5.26 $Y=0.79
c104 23 0 1.14729e-19 $X=4.905 $Y=2.08
c105 4 0 1.47738e-19 $X=5.355 $Y=2.155
r106 35 38 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.99 $Y=0.79
+ $X2=5.26 $Y2=0.79
r107 29 31 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.075 $Y=2.605
+ $X2=5.495 $Y2=2.605
r108 28 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.99 $Y=2.44
+ $X2=5.075 $Y2=2.605
r109 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=2.165
+ $X2=4.99 $Y2=2.08
r110 27 28 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.99 $Y=2.165
+ $X2=4.99 $Y2=2.44
r111 26 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=1.995
+ $X2=4.99 $Y2=2.08
r112 25 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=0.955
+ $X2=4.99 $Y2=0.79
r113 25 26 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.99 $Y=0.955
+ $X2=4.99 $Y2=1.995
r114 23 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=2.08
+ $X2=4.99 $Y2=2.08
r115 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.905 $Y=2.08
+ $X2=4.215 $Y2=2.08
r116 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.13 $Y=2.165
+ $X2=4.215 $Y2=2.08
r117 21 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.13 $Y=2.165
+ $X2=4.13 $Y2=2.37
r118 20 34 3.6737 $w=1.7e-07 $l=1.33604e-07 $layer=LI1_cond $X=1.245 $Y=2.455
+ $X2=1.14 $Y2=2.52
r119 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.045 $Y=2.455
+ $X2=4.13 $Y2=2.37
r120 19 20 182.674 $w=1.68e-07 $l=2.8e-06 $layer=LI1_cond $X=4.045 $Y=2.455
+ $X2=1.245 $Y2=2.455
r121 15 18 71.8268 $w=2.08e-07 $l=1.36e-06 $layer=LI1_cond $X=1.14 $Y=0.805
+ $X2=1.14 $Y2=2.165
r122 13 34 3.2415 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=1.14 $Y=2.37 $X2=1.14
+ $Y2=2.52
r123 13 18 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=1.14 $Y=2.37
+ $X2=1.14 $Y2=2.165
r124 4 31 600 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=2.155 $X2=5.495 $Y2=2.605
r125 3 34 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=2.01 $X2=1.14 $Y2=2.505
r126 3 18 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=2.01 $X2=1.14 $Y2=2.165
r127 2 38 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=5.12
+ $Y=0.595 $X2=5.26 $Y2=0.79
r128 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.595 $X2=1.14 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 45 57 61 77 78 81 84
r103 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r104 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r105 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r106 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r107 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r108 72 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r109 72 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 71 74 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r111 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r112 69 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.435 $Y2=3.33
r113 69 71 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 68 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r115 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r116 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r117 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r118 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 62 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 61 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.27 $Y=3.33
+ $X2=6.435 $Y2=3.33
r122 61 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.27 $Y=3.33 $X2=6
+ $Y2=3.33
r123 60 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r124 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 57 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 57 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.395 $Y=3.33
+ $X2=4.08 $Y2=3.33
r127 56 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r128 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r129 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r130 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r131 49 53 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r132 48 52 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r133 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r134 45 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r135 45 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 43 74 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.49 $Y=3.33 $X2=8.4
+ $Y2=3.33
r137 43 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.49 $Y=3.33
+ $X2=8.595 $Y2=3.33
r138 42 77 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.7 $Y=3.33
+ $X2=9.36 $Y2=3.33
r139 42 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.7 $Y=3.33
+ $X2=8.595 $Y2=3.33
r140 40 55 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.12 $Y2=3.33
r141 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.35 $Y2=3.33
r142 39 59 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.35 $Y2=3.33
r144 37 52 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.49 $Y2=3.33
r146 36 55 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=3.12 $Y2=3.33
r147 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=2.49 $Y2=3.33
r148 32 44 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.595 $Y=3.245
+ $X2=8.595 $Y2=3.33
r149 32 34 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=8.595 $Y=3.245
+ $X2=8.595 $Y2=2.59
r150 28 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=3.245
+ $X2=6.435 $Y2=3.33
r151 28 30 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=6.435 $Y=3.245
+ $X2=6.435 $Y2=2.59
r152 24 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.56 $Y2=3.33
r153 24 26 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.56 $Y2=2.45
r154 20 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=3.245
+ $X2=3.35 $Y2=3.33
r155 20 22 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.35 $Y=3.245
+ $X2=3.35 $Y2=2.81
r156 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=3.33
r157 16 18 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=2.81
r158 5 34 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=8.455
+ $Y=2.095 $X2=8.595 $Y2=2.59
r159 4 30 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=2.095 $X2=6.435 $Y2=2.59
r160 3 26 300 $w=1.7e-07 $l=9.90139e-07 $layer=licon1_PDIFF $count=2 $X=4.07
+ $Y=1.675 $X2=4.56 $Y2=2.45
r161 2 22 600 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.675 $X2=3.35 $Y2=2.81
r162 1 18 600 $w=1.7e-07 $l=1.25605e-06 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.675 $X2=2.49 $Y2=2.81
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%X 1 2 3 4 13 19 21 22 25 29 30 37 45
c54 29 0 2.62564e-19 $X=3.995 $Y=1.21
r55 36 45 2.49696 $w=2.98e-07 $l=6.5e-08 $layer=LI1_cond $X=4.015 $Y=1.36
+ $X2=4.015 $Y2=1.295
r56 30 37 3.56541 $w=3e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.93 $Y=1.815
+ $X2=4.015 $Y2=1.645
r57 30 37 1.26769 $w=2.98e-07 $l=3.3e-08 $layer=LI1_cond $X=4.015 $Y=1.612
+ $X2=4.015 $Y2=1.645
r58 29 45 0.384148 $w=2.98e-07 $l=1e-08 $layer=LI1_cond $X=4.015 $Y=1.285
+ $X2=4.015 $Y2=1.295
r59 29 30 9.29637 $w=2.98e-07 $l=2.42e-07 $layer=LI1_cond $X=4.015 $Y=1.37
+ $X2=4.015 $Y2=1.612
r60 29 36 0.384148 $w=2.98e-07 $l=1e-08 $layer=LI1_cond $X=4.015 $Y=1.37
+ $X2=4.015 $Y2=1.36
r61 27 29 9.94137 $w=2.08e-07 $l=1.8e-07 $layer=LI1_cond $X=3.95 $Y=1.03
+ $X2=3.95 $Y2=1.21
r62 27 28 4.70473 $w=1.9e-07 $l=9.44722e-08 $layer=LI1_cond $X=3.95 $Y=1.03
+ $X2=3.93 $Y2=0.945
r63 23 28 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=0.86 $X2=3.93
+ $Y2=0.945
r64 23 25 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.93 $Y=0.86
+ $X2=3.93 $Y2=0.525
r65 21 28 1.74598 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.825 $Y=0.945
+ $X2=3.93 $Y2=0.945
r66 21 22 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.825 $Y=0.945
+ $X2=3.175 $Y2=0.945
r67 17 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.07 $Y=0.86
+ $X2=3.175 $Y2=0.945
r68 17 19 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.07 $Y=0.86
+ $X2=3.07 $Y2=0.525
r69 13 30 3.28577 $w=3.4e-07 $l=2.35e-07 $layer=LI1_cond $X=3.695 $Y=1.815
+ $X2=3.93 $Y2=1.815
r70 13 15 26.2689 $w=3.38e-07 $l=7.75e-07 $layer=LI1_cond $X=3.695 $Y=1.815
+ $X2=2.92 $Y2=1.815
r71 4 30 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.64
+ $Y=1.675 $X2=3.78 $Y2=1.82
r72 3 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.675 $X2=2.92 $Y2=1.82
r73 2 25 91 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=2 $X=3.79
+ $Y=0.235 $X2=3.93 $Y2=0.525
r74 1 19 91 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=2 $X=2.93
+ $Y=0.235 $X2=3.07 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 45 47 62 77 78 81 84
r119 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r120 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r121 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r122 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r123 74 77 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r124 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r125 72 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r126 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r127 69 72 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r128 69 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r129 68 71 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r130 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r131 66 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.13
+ $Y2=0
r132 66 68 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.295 $Y=0
+ $X2=6.48 $Y2=0
r133 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r134 62 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=0 $X2=6.13
+ $Y2=0
r135 62 64 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=4.56 $Y2=0
r136 61 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r137 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r138 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r139 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r140 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r141 55 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.65
+ $Y2=0
r142 55 57 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.12 $Y2=0
r143 54 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r144 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r145 50 54 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=2.16 $Y2=0
r146 49 53 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r147 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r148 47 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.555 $Y=0 $X2=2.65
+ $Y2=0
r149 47 53 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=0
+ $X2=2.16 $Y2=0
r150 45 85 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=6
+ $Y2=0
r151 45 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r152 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=0 $X2=8.4
+ $Y2=0
r153 43 71 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=7.92
+ $Y2=0
r154 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.235
+ $Y2=0
r155 40 60 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.255 $Y=0
+ $X2=4.08 $Y2=0
r156 40 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.36
+ $Y2=0
r157 39 64 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.56
+ $Y2=0
r158 39 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.36
+ $Y2=0
r159 37 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=0
+ $X2=3.12 $Y2=0
r160 37 38 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.5
+ $Y2=0
r161 36 60 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=0
+ $X2=4.08 $Y2=0
r162 36 38 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.605 $Y=0 $X2=3.5
+ $Y2=0
r163 32 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.235 $Y=0.085
+ $X2=8.235 $Y2=0
r164 32 34 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=8.235 $Y=0.085
+ $X2=8.235 $Y2=0.74
r165 28 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0
r166 28 30 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0.615
r167 24 41 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.36 $Y=0.085
+ $X2=4.36 $Y2=0
r168 24 26 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.36 $Y=0.085
+ $X2=4.36 $Y2=0.38
r169 20 38 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=0.085
+ $X2=3.5 $Y2=0
r170 20 22 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.5 $Y=0.085
+ $X2=3.5 $Y2=0.38
r171 16 81 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0
r172 16 18 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.65 $Y=0.085
+ $X2=2.65 $Y2=0.38
r173 5 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.095
+ $Y=0.595 $X2=8.235 $Y2=0.74
r174 4 30 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.595 $X2=6.13 $Y2=0.615
r175 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.22
+ $Y=0.235 $X2=4.36 $Y2=0.38
r176 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.36
+ $Y=0.235 $X2=3.5 $Y2=0.38
r177 1 18 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.655 $X2=2.64 $Y2=0.38
.ends

