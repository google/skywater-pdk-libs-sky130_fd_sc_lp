* File: sky130_fd_sc_lp__and4b_m.pxi.spice
* Created: Fri Aug 28 10:08:56 2020
* 
x_PM_SKY130_FD_SC_LP__AND4B_M%A_N N_A_N_M1007_g N_A_N_c_84_n N_A_N_c_85_n
+ N_A_N_c_86_n N_A_N_M1008_g N_A_N_c_81_n A_N N_A_N_c_82_n N_A_N_c_83_n
+ PM_SKY130_FD_SC_LP__AND4B_M%A_N
x_PM_SKY130_FD_SC_LP__AND4B_M%A_27_55# N_A_27_55#_M1007_s N_A_27_55#_M1008_s
+ N_A_27_55#_c_119_n N_A_27_55#_c_120_n N_A_27_55#_c_121_n N_A_27_55#_c_122_n
+ N_A_27_55#_c_123_n N_A_27_55#_c_133_n N_A_27_55#_M1010_g N_A_27_55#_c_124_n
+ N_A_27_55#_M1002_g N_A_27_55#_c_125_n N_A_27_55#_c_126_n N_A_27_55#_c_134_n
+ N_A_27_55#_c_127_n N_A_27_55#_c_128_n N_A_27_55#_c_129_n N_A_27_55#_c_135_n
+ N_A_27_55#_c_130_n N_A_27_55#_c_131_n N_A_27_55#_c_137_n
+ PM_SKY130_FD_SC_LP__AND4B_M%A_27_55#
x_PM_SKY130_FD_SC_LP__AND4B_M%B N_B_M1003_g N_B_M1001_g B B B N_B_c_201_n
+ PM_SKY130_FD_SC_LP__AND4B_M%B
x_PM_SKY130_FD_SC_LP__AND4B_M%C N_C_M1004_g N_C_M1005_g N_C_c_233_n N_C_c_234_n
+ N_C_c_235_n C C C N_C_c_237_n PM_SKY130_FD_SC_LP__AND4B_M%C
x_PM_SKY130_FD_SC_LP__AND4B_M%D N_D_M1009_g N_D_M1006_g N_D_c_271_n N_D_c_272_n
+ N_D_c_273_n D D N_D_c_275_n PM_SKY130_FD_SC_LP__AND4B_M%D
x_PM_SKY130_FD_SC_LP__AND4B_M%A_240_73# N_A_240_73#_M1002_s N_A_240_73#_M1010_d
+ N_A_240_73#_M1005_d N_A_240_73#_c_306_n N_A_240_73#_M1011_g
+ N_A_240_73#_M1000_g N_A_240_73#_c_305_n N_A_240_73#_c_309_n
+ N_A_240_73#_c_310_n N_A_240_73#_c_311_n N_A_240_73#_c_312_n
+ N_A_240_73#_c_313_n N_A_240_73#_c_314_n PM_SKY130_FD_SC_LP__AND4B_M%A_240_73#
x_PM_SKY130_FD_SC_LP__AND4B_M%VPWR N_VPWR_M1008_d N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n
+ VPWR N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_375_n
+ N_VPWR_c_385_n N_VPWR_c_386_n PM_SKY130_FD_SC_LP__AND4B_M%VPWR
x_PM_SKY130_FD_SC_LP__AND4B_M%X N_X_M1011_d N_X_M1000_d X X X X X X X
+ PM_SKY130_FD_SC_LP__AND4B_M%X
x_PM_SKY130_FD_SC_LP__AND4B_M%VGND N_VGND_M1007_d N_VGND_M1009_d N_VGND_c_430_n
+ N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n VGND N_VGND_c_434_n
+ N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n PM_SKY130_FD_SC_LP__AND4B_M%VGND
cc_1 VNB N_A_N_M1007_g 0.0324801f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.485
cc_2 VNB N_A_N_c_81_n 0.0430651f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.715
cc_3 VNB N_A_N_c_82_n 0.0190717f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_4 VNB N_A_N_c_83_n 0.0266584f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_5 VNB N_A_27_55#_c_119_n 0.0362426f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.195
cc_6 VNB N_A_27_55#_c_120_n 0.0108611f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_7 VNB N_A_27_55#_c_121_n 0.0270057f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.975
cc_8 VNB N_A_27_55#_c_122_n 0.0132586f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.715
cc_9 VNB N_A_27_55#_c_123_n 0.0120437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_55#_c_124_n 0.0204864f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.31
cc_11 VNB N_A_27_55#_c_125_n 0.0302562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_55#_c_126_n 0.0248172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_55#_c_127_n 4.08405e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_55#_c_128_n 0.0121159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_55#_c_129_n 0.00869196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_55#_c_130_n 0.00286107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_55#_c_131_n 0.0167702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_M1003_g 0.0313132f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.485
cc_19 VNB N_B_M1001_g 0.00961741f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.865
cc_20 VNB B 0.00675676f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.195
cc_21 VNB N_B_c_201_n 0.033218f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_22 VNB N_C_M1005_g 0.00496318f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.79
cc_23 VNB N_C_c_233_n 0.0168693f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.195
cc_24 VNB N_C_c_234_n 0.0209027f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_25 VNB N_C_c_235_n 0.0151455f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.975
cc_26 VNB C 0.00809908f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.715
cc_27 VNB N_C_c_237_n 0.0174736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_D_M1006_g 0.00525575f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.79
cc_29 VNB N_D_c_271_n 0.0185981f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.195
cc_30 VNB N_D_c_272_n 0.0209027f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_31 VNB N_D_c_273_n 0.0153418f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.975
cc_32 VNB D 0.0164107f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.715
cc_33 VNB N_D_c_275_n 0.0153418f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_34 VNB N_A_240_73#_M1011_g 0.0637345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_240_73#_c_305_n 0.0111197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_375_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB X 0.0559917f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.865
cc_38 VNB N_VGND_c_430_n 0.00696239f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.195
cc_39 VNB N_VGND_c_431_n 0.00643792f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_40 VNB N_VGND_c_432_n 0.0574372f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_41 VNB N_VGND_c_433_n 0.00609509f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.14
cc_42 VNB N_VGND_c_434_n 0.0159906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_435_n 0.021708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_436_n 0.241049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_437_n 0.00540805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_A_N_c_84_n 0.0382998f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.79
cc_47 VPB N_A_N_c_85_n 0.0317838f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.79
cc_48 VPB N_A_N_c_86_n 0.024167f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.865
cc_49 VPB N_A_N_c_81_n 0.00662274f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.715
cc_50 VPB N_A_27_55#_c_123_n 0.00450173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_27_55#_c_133_n 0.0190554f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.14
cc_52 VPB N_A_27_55#_c_134_n 0.0160698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_55#_c_135_n 0.00349719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_27_55#_c_130_n 0.00104057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_27_55#_c_137_n 0.00365811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_B_M1001_g 0.0289393f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.865
cc_57 VPB N_C_M1005_g 0.0288696f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.79
cc_58 VPB N_D_M1006_g 0.0296913f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.79
cc_59 VPB N_A_240_73#_c_306_n 0.0472251f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.14
cc_60 VPB N_A_240_73#_M1011_g 0.0415614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_240_73#_c_305_n 8.70082e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_240_73#_c_309_n 0.00179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_240_73#_c_310_n 0.0223695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_240_73#_c_311_n 0.00982935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_240_73#_c_312_n 0.00255537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_240_73#_c_313_n 0.00912535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_240_73#_c_314_n 0.0461649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_376_n 0.0397419f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.715
cc_69 VPB N_VPWR_c_377_n 0.0225617f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.14
cc_70 VPB N_VPWR_c_378_n 0.019582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_379_n 0.0193975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_380_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_381_n 0.0374657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_382_n 0.0203024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_383_n 0.0210716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_375_n 0.119996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_385_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_386_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.0584189f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.865
cc_80 N_A_N_M1007_g N_A_27_55#_c_120_n 0.0136976f $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_81 N_A_N_c_84_n N_A_27_55#_c_122_n 0.0188644f $X=0.925 $Y=1.79 $X2=0 $Y2=0
cc_82 N_A_N_c_81_n N_A_27_55#_c_122_n 0.0145557f $X=0.385 $Y=1.715 $X2=0 $Y2=0
cc_83 N_A_N_c_84_n N_A_27_55#_c_123_n 0.00521434f $X=0.925 $Y=1.79 $X2=0 $Y2=0
cc_84 N_A_N_c_86_n N_A_27_55#_c_133_n 0.0108557f $X=1 $Y=1.865 $X2=0 $Y2=0
cc_85 N_A_N_c_82_n N_A_27_55#_c_126_n 0.0145557f $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_86 N_A_N_c_83_n N_A_27_55#_c_126_n 0.00167181f $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_87 N_A_N_c_86_n N_A_27_55#_c_134_n 0.00521434f $X=1 $Y=1.865 $X2=0 $Y2=0
cc_88 N_A_N_M1007_g N_A_27_55#_c_127_n 3.52891e-19 $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_89 N_A_N_M1007_g N_A_27_55#_c_128_n 0.013224f $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_90 N_A_N_c_82_n N_A_27_55#_c_128_n 0.00157812f $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_91 N_A_N_c_83_n N_A_27_55#_c_128_n 0.0146605f $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_92 N_A_N_c_82_n N_A_27_55#_c_129_n 0.00368742f $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_93 N_A_N_c_83_n N_A_27_55#_c_129_n 0.0157003f $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_94 N_A_N_c_84_n N_A_27_55#_c_135_n 0.00196805f $X=0.925 $Y=1.79 $X2=0 $Y2=0
cc_95 N_A_N_c_86_n N_A_27_55#_c_135_n 0.00282651f $X=1 $Y=1.865 $X2=0 $Y2=0
cc_96 N_A_N_M1007_g N_A_27_55#_c_130_n 0.00103261f $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_97 N_A_N_c_84_n N_A_27_55#_c_130_n 0.00420973f $X=0.925 $Y=1.79 $X2=0 $Y2=0
cc_98 N_A_N_c_81_n N_A_27_55#_c_130_n 0.00553214f $X=0.385 $Y=1.715 $X2=0 $Y2=0
cc_99 N_A_N_c_82_n N_A_27_55#_c_130_n 4.73066e-19 $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_100 N_A_N_c_83_n N_A_27_55#_c_130_n 0.0243898f $X=0.385 $Y=1.14 $X2=0 $Y2=0
cc_101 N_A_N_M1007_g N_A_27_55#_c_131_n 0.0145557f $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_102 N_A_N_c_84_n N_A_27_55#_c_137_n 0.0179614f $X=0.925 $Y=1.79 $X2=0 $Y2=0
cc_103 N_A_N_c_86_n N_A_27_55#_c_137_n 0.00527066f $X=1 $Y=1.865 $X2=0 $Y2=0
cc_104 N_A_N_c_84_n N_A_240_73#_c_305_n 2.02157e-19 $X=0.925 $Y=1.79 $X2=0 $Y2=0
cc_105 N_A_N_c_84_n N_A_240_73#_c_311_n 0.00128646f $X=0.925 $Y=1.79 $X2=0 $Y2=0
cc_106 N_A_N_c_86_n N_VPWR_c_376_n 0.003345f $X=1 $Y=1.865 $X2=0 $Y2=0
cc_107 N_A_N_c_86_n N_VPWR_c_375_n 0.00393927f $X=1 $Y=1.865 $X2=0 $Y2=0
cc_108 N_A_N_M1007_g N_VGND_c_430_n 0.0121979f $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_109 N_A_N_M1007_g N_VGND_c_434_n 0.00334249f $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_110 N_A_N_M1007_g N_VGND_c_436_n 0.00484861f $X=0.475 $Y=0.485 $X2=0 $Y2=0
cc_111 N_A_27_55#_c_119_n N_B_M1003_g 0.0442408f $X=1.465 $Y=0.18 $X2=0 $Y2=0
cc_112 N_A_27_55#_c_123_n N_B_M1001_g 0.00723725f $X=1.36 $Y=1.725 $X2=0 $Y2=0
cc_113 N_A_27_55#_c_134_n N_B_M1001_g 0.0189045f $X=1.46 $Y=1.8 $X2=0 $Y2=0
cc_114 N_A_27_55#_c_121_n B 0.00101947f $X=1.285 $Y=1.4 $X2=0 $Y2=0
cc_115 N_A_27_55#_c_124_n B 0.0094098f $X=1.54 $Y=0.255 $X2=0 $Y2=0
cc_116 N_A_27_55#_c_121_n N_B_c_201_n 0.010441f $X=1.285 $Y=1.4 $X2=0 $Y2=0
cc_117 N_A_27_55#_c_126_n N_B_c_201_n 0.00119702f $X=0.925 $Y=1.325 $X2=0 $Y2=0
cc_118 N_A_27_55#_c_119_n N_A_240_73#_c_305_n 0.00336639f $X=1.465 $Y=0.18 $X2=0
+ $Y2=0
cc_119 N_A_27_55#_c_121_n N_A_240_73#_c_305_n 0.0115398f $X=1.285 $Y=1.4 $X2=0
+ $Y2=0
cc_120 N_A_27_55#_c_123_n N_A_240_73#_c_305_n 0.010194f $X=1.36 $Y=1.725 $X2=0
+ $Y2=0
cc_121 N_A_27_55#_c_124_n N_A_240_73#_c_305_n 0.00110123f $X=1.54 $Y=0.255 $X2=0
+ $Y2=0
cc_122 N_A_27_55#_c_125_n N_A_240_73#_c_305_n 0.0129654f $X=0.925 $Y=0.805 $X2=0
+ $Y2=0
cc_123 N_A_27_55#_c_134_n N_A_240_73#_c_305_n 9.9455e-19 $X=1.46 $Y=1.8 $X2=0
+ $Y2=0
cc_124 N_A_27_55#_c_128_n N_A_240_73#_c_305_n 0.0115207f $X=0.84 $Y=0.79 $X2=0
+ $Y2=0
cc_125 N_A_27_55#_c_130_n N_A_240_73#_c_305_n 0.0538665f $X=0.925 $Y=0.97 $X2=0
+ $Y2=0
cc_126 N_A_27_55#_c_133_n N_A_240_73#_c_309_n 0.00177249f $X=1.46 $Y=1.875 $X2=0
+ $Y2=0
cc_127 N_A_27_55#_c_121_n N_A_240_73#_c_311_n 2.35045e-19 $X=1.285 $Y=1.4 $X2=0
+ $Y2=0
cc_128 N_A_27_55#_c_133_n N_A_240_73#_c_311_n 0.00770346f $X=1.46 $Y=1.875 $X2=0
+ $Y2=0
cc_129 N_A_27_55#_c_134_n N_A_240_73#_c_311_n 0.0116323f $X=1.46 $Y=1.8 $X2=0
+ $Y2=0
cc_130 N_A_27_55#_c_137_n N_A_240_73#_c_311_n 0.0121076f $X=0.925 $Y=1.83 $X2=0
+ $Y2=0
cc_131 N_A_27_55#_c_121_n N_VPWR_c_376_n 0.00250436f $X=1.285 $Y=1.4 $X2=0 $Y2=0
cc_132 N_A_27_55#_c_133_n N_VPWR_c_376_n 0.003503f $X=1.46 $Y=1.875 $X2=0 $Y2=0
cc_133 N_A_27_55#_c_134_n N_VPWR_c_376_n 2.39228e-19 $X=1.46 $Y=1.8 $X2=0 $Y2=0
cc_134 N_A_27_55#_c_133_n N_VPWR_c_377_n 7.00463e-19 $X=1.46 $Y=1.875 $X2=0
+ $Y2=0
cc_135 N_A_27_55#_c_133_n N_VPWR_c_375_n 0.00393928f $X=1.46 $Y=1.875 $X2=0
+ $Y2=0
cc_136 N_A_27_55#_c_120_n N_VGND_c_430_n 0.0107746f $X=1.09 $Y=0.18 $X2=0 $Y2=0
cc_137 N_A_27_55#_c_128_n N_VGND_c_430_n 0.022235f $X=0.84 $Y=0.79 $X2=0 $Y2=0
cc_138 N_A_27_55#_c_131_n N_VGND_c_430_n 5.81838e-19 $X=0.925 $Y=0.97 $X2=0
+ $Y2=0
cc_139 N_A_27_55#_c_120_n N_VGND_c_432_n 0.0223042f $X=1.09 $Y=0.18 $X2=0 $Y2=0
cc_140 N_A_27_55#_c_128_n N_VGND_c_432_n 0.00256533f $X=0.84 $Y=0.79 $X2=0 $Y2=0
cc_141 N_A_27_55#_c_127_n N_VGND_c_434_n 0.00696263f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_142 N_A_27_55#_c_128_n N_VGND_c_434_n 0.00259759f $X=0.84 $Y=0.79 $X2=0 $Y2=0
cc_143 N_A_27_55#_c_119_n N_VGND_c_436_n 0.0266423f $X=1.465 $Y=0.18 $X2=0 $Y2=0
cc_144 N_A_27_55#_c_120_n N_VGND_c_436_n 0.00849369f $X=1.09 $Y=0.18 $X2=0 $Y2=0
cc_145 N_A_27_55#_c_127_n N_VGND_c_436_n 0.00670996f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_146 N_A_27_55#_c_128_n N_VGND_c_436_n 0.00975009f $X=0.84 $Y=0.79 $X2=0 $Y2=0
cc_147 N_B_M1001_g N_C_M1005_g 0.0272599f $X=1.9 $Y=2.195 $X2=0 $Y2=0
cc_148 N_B_M1003_g N_C_c_233_n 0.0268594f $X=1.9 $Y=0.575 $X2=0 $Y2=0
cc_149 B N_C_c_233_n 9.11751e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_150 N_B_M1001_g N_C_c_234_n 0.0268594f $X=1.9 $Y=2.195 $X2=0 $Y2=0
cc_151 N_B_M1003_g C 0.00741039f $X=1.9 $Y=0.575 $X2=0 $Y2=0
cc_152 B C 0.0764259f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_153 N_B_c_201_n N_C_c_237_n 0.0268594f $X=1.81 $Y=1.32 $X2=0 $Y2=0
cc_154 N_B_M1003_g N_A_240_73#_c_305_n 0.001167f $X=1.9 $Y=0.575 $X2=0 $Y2=0
cc_155 N_B_M1001_g N_A_240_73#_c_305_n 0.00128518f $X=1.9 $Y=2.195 $X2=0 $Y2=0
cc_156 B N_A_240_73#_c_305_n 0.0618037f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_157 N_B_c_201_n N_A_240_73#_c_305_n 0.00100646f $X=1.81 $Y=1.32 $X2=0 $Y2=0
cc_158 N_B_M1001_g N_A_240_73#_c_309_n 0.00174999f $X=1.9 $Y=2.195 $X2=0 $Y2=0
cc_159 N_B_M1001_g N_A_240_73#_c_310_n 0.0172266f $X=1.9 $Y=2.195 $X2=0 $Y2=0
cc_160 B N_A_240_73#_c_311_n 0.0172269f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_161 N_B_c_201_n N_A_240_73#_c_311_n 0.00115776f $X=1.81 $Y=1.32 $X2=0 $Y2=0
cc_162 N_B_M1001_g N_VPWR_c_377_n 0.00795896f $X=1.9 $Y=2.195 $X2=0 $Y2=0
cc_163 N_B_M1001_g N_VPWR_c_375_n 0.00357161f $X=1.9 $Y=2.195 $X2=0 $Y2=0
cc_164 N_B_M1003_g N_VGND_c_432_n 0.00393992f $X=1.9 $Y=0.575 $X2=0 $Y2=0
cc_165 B N_VGND_c_432_n 0.0069537f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_166 N_B_M1003_g N_VGND_c_436_n 0.0067116f $X=1.9 $Y=0.575 $X2=0 $Y2=0
cc_167 B N_VGND_c_436_n 0.00973813f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_168 B A_323_73# 0.00139886f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_169 N_C_M1005_g N_D_M1006_g 0.0231099f $X=2.345 $Y=2.195 $X2=0 $Y2=0
cc_170 N_C_c_233_n N_D_c_271_n 0.0187918f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_171 C N_D_c_271_n 0.00648897f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_172 N_C_c_234_n N_D_c_272_n 0.013969f $X=2.35 $Y=1.4 $X2=0 $Y2=0
cc_173 N_C_c_235_n N_D_c_273_n 0.013969f $X=2.35 $Y=1.565 $X2=0 $Y2=0
cc_174 C D 0.0298848f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_175 N_C_c_237_n D 0.00216519f $X=2.35 $Y=1.06 $X2=0 $Y2=0
cc_176 C N_D_c_275_n 0.0021666f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_177 N_C_c_237_n N_D_c_275_n 0.013969f $X=2.35 $Y=1.06 $X2=0 $Y2=0
cc_178 C N_A_240_73#_c_305_n 0.00215796f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_179 N_C_M1005_g N_A_240_73#_c_310_n 0.0141804f $X=2.345 $Y=2.195 $X2=0 $Y2=0
cc_180 N_C_c_235_n N_A_240_73#_c_310_n 0.00419575f $X=2.35 $Y=1.565 $X2=0 $Y2=0
cc_181 C N_A_240_73#_c_310_n 0.0273269f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_182 N_C_M1005_g N_A_240_73#_c_313_n 0.00737656f $X=2.345 $Y=2.195 $X2=0 $Y2=0
cc_183 N_C_M1005_g N_VPWR_c_377_n 0.00627777f $X=2.345 $Y=2.195 $X2=0 $Y2=0
cc_184 N_C_M1005_g N_VPWR_c_375_n 0.0034403f $X=2.345 $Y=2.195 $X2=0 $Y2=0
cc_185 N_C_c_233_n N_VGND_c_431_n 0.00124648f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_186 C N_VGND_c_431_n 0.00569849f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_187 N_C_c_233_n N_VGND_c_432_n 0.00309992f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_188 C N_VGND_c_432_n 0.00859527f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_189 N_C_c_233_n N_VGND_c_436_n 0.00387028f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_190 C N_VGND_c_436_n 0.0114764f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_191 C A_395_73# 0.00345969f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_192 C A_467_73# 0.00488434f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_193 N_D_M1006_g N_A_240_73#_M1011_g 0.0215315f $X=2.8 $Y=2.195 $X2=0 $Y2=0
cc_194 N_D_c_271_n N_A_240_73#_M1011_g 0.0135161f $X=2.89 $Y=0.895 $X2=0 $Y2=0
cc_195 D N_A_240_73#_M1011_g 0.00583598f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_196 N_D_c_275_n N_A_240_73#_M1011_g 0.0391028f $X=2.89 $Y=1.06 $X2=0 $Y2=0
cc_197 N_D_M1006_g N_A_240_73#_c_310_n 0.00557179f $X=2.8 $Y=2.195 $X2=0 $Y2=0
cc_198 N_D_M1006_g N_A_240_73#_c_312_n 5.45931e-19 $X=2.8 $Y=2.195 $X2=0 $Y2=0
cc_199 N_D_M1006_g N_A_240_73#_c_313_n 0.00340996f $X=2.8 $Y=2.195 $X2=0 $Y2=0
cc_200 N_D_M1006_g N_A_240_73#_c_314_n 0.00953828f $X=2.8 $Y=2.195 $X2=0 $Y2=0
cc_201 N_D_M1006_g N_VPWR_c_378_n 0.00407252f $X=2.8 $Y=2.195 $X2=0 $Y2=0
cc_202 N_D_c_273_n N_VPWR_c_378_n 4.18433e-19 $X=2.89 $Y=1.565 $X2=0 $Y2=0
cc_203 D N_VPWR_c_378_n 0.00811988f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_204 D X 0.0462346f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_205 N_D_c_271_n N_VGND_c_431_n 0.00952047f $X=2.89 $Y=0.895 $X2=0 $Y2=0
cc_206 D N_VGND_c_431_n 0.0210792f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_207 N_D_c_275_n N_VGND_c_431_n 0.00101918f $X=2.89 $Y=1.06 $X2=0 $Y2=0
cc_208 N_D_c_271_n N_VGND_c_432_n 0.00386543f $X=2.89 $Y=0.895 $X2=0 $Y2=0
cc_209 N_D_c_271_n N_VGND_c_436_n 0.00629974f $X=2.89 $Y=0.895 $X2=0 $Y2=0
cc_210 D N_VGND_c_436_n 0.00377899f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_211 N_A_240_73#_c_311_n N_VPWR_c_376_n 0.00781527f $X=1.78 $Y=1.83 $X2=0
+ $Y2=0
cc_212 N_A_240_73#_c_310_n N_VPWR_c_377_n 0.0168901f $X=2.48 $Y=1.83 $X2=0 $Y2=0
cc_213 N_A_240_73#_c_312_n N_VPWR_c_377_n 0.0122852f $X=2.585 $Y=2.855 $X2=0
+ $Y2=0
cc_214 N_A_240_73#_c_313_n N_VPWR_c_377_n 0.0498507f $X=2.585 $Y=2.13 $X2=0
+ $Y2=0
cc_215 N_A_240_73#_c_314_n N_VPWR_c_377_n 0.00635329f $X=2.645 $Y=2.85 $X2=0
+ $Y2=0
cc_216 N_A_240_73#_c_306_n N_VPWR_c_378_n 0.0186987f $X=3.265 $Y=2.85 $X2=0
+ $Y2=0
cc_217 N_A_240_73#_M1011_g N_VPWR_c_378_n 0.00799165f $X=3.34 $Y=0.575 $X2=0
+ $Y2=0
cc_218 N_A_240_73#_c_312_n N_VPWR_c_378_n 0.0120815f $X=2.585 $Y=2.855 $X2=0
+ $Y2=0
cc_219 N_A_240_73#_c_313_n N_VPWR_c_378_n 0.0305673f $X=2.585 $Y=2.13 $X2=0
+ $Y2=0
cc_220 N_A_240_73#_c_314_n N_VPWR_c_378_n 0.00358618f $X=2.645 $Y=2.85 $X2=0
+ $Y2=0
cc_221 N_A_240_73#_c_306_n N_VPWR_c_379_n 0.00445258f $X=3.265 $Y=2.85 $X2=0
+ $Y2=0
cc_222 N_A_240_73#_c_312_n N_VPWR_c_379_n 0.0152941f $X=2.585 $Y=2.855 $X2=0
+ $Y2=0
cc_223 N_A_240_73#_c_314_n N_VPWR_c_379_n 0.00593936f $X=2.645 $Y=2.85 $X2=0
+ $Y2=0
cc_224 N_A_240_73#_c_306_n N_VPWR_c_383_n 0.00625242f $X=3.265 $Y=2.85 $X2=0
+ $Y2=0
cc_225 N_A_240_73#_c_306_n N_VPWR_c_375_n 0.0114224f $X=3.265 $Y=2.85 $X2=0
+ $Y2=0
cc_226 N_A_240_73#_c_312_n N_VPWR_c_375_n 0.0104794f $X=2.585 $Y=2.855 $X2=0
+ $Y2=0
cc_227 N_A_240_73#_c_314_n N_VPWR_c_375_n 0.00814482f $X=2.645 $Y=2.85 $X2=0
+ $Y2=0
cc_228 N_A_240_73#_M1011_g X 0.0500664f $X=3.34 $Y=0.575 $X2=0 $Y2=0
cc_229 N_A_240_73#_c_305_n N_VGND_c_430_n 0.00227392f $X=1.325 $Y=0.64 $X2=0
+ $Y2=0
cc_230 N_A_240_73#_M1011_g N_VGND_c_431_n 0.0078198f $X=3.34 $Y=0.575 $X2=0
+ $Y2=0
cc_231 N_A_240_73#_c_305_n N_VGND_c_432_n 0.00534682f $X=1.325 $Y=0.64 $X2=0
+ $Y2=0
cc_232 N_A_240_73#_M1011_g N_VGND_c_435_n 0.00465548f $X=3.34 $Y=0.575 $X2=0
+ $Y2=0
cc_233 N_A_240_73#_M1011_g N_VGND_c_436_n 0.00927152f $X=3.34 $Y=0.575 $X2=0
+ $Y2=0
cc_234 N_A_240_73#_c_305_n N_VGND_c_436_n 0.00564111f $X=1.325 $Y=0.64 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_378_n X 0.0356067f $X=3.095 $Y=2.26 $X2=0 $Y2=0
cc_236 N_VPWR_c_383_n X 0.00698589f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_237 N_VPWR_c_375_n X 0.00795962f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_238 X N_VGND_c_435_n 0.00646233f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_239 X N_VGND_c_436_n 0.00795962f $X=3.515 $Y=0.47 $X2=0 $Y2=0
