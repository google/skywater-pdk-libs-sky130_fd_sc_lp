* File: sky130_fd_sc_lp__sleep_pargate_plv_21.pxi.spice
* Created: Wed Sep  2 10:37:41 2020
* 
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%SLEEP N_SLEEP_c_38_n N_SLEEP_M1000_g
+ N_SLEEP_c_39_n N_SLEEP_M1001_g N_SLEEP_c_40_n N_SLEEP_M1002_g N_SLEEP_c_41_n
+ SLEEP SLEEP SLEEP SLEEP SLEEP N_SLEEP_c_43_n N_SLEEP_c_44_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%SLEEP
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%VPWR N_VPWR_M1000_s N_VPWR_M1001_s
+ VPWR N_VPWR_c_93_n N_VPWR_c_94_n N_VPWR_c_95_n N_VPWR_c_96_n N_VPWR_c_97_n
+ N_VPWR_c_98_n N_VPWR_c_99_n N_VPWR_c_92_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%VPWR
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%VIRTPWR N_VIRTPWR_M1000_d
+ N_VIRTPWR_M1002_d N_VIRTPWR_c_190_n N_VIRTPWR_c_191_n VIRTPWR
+ N_VIRTPWR_c_192_n N_VIRTPWR_c_193_n N_VIRTPWR_c_194_n N_VIRTPWR_c_195_n
+ N_VIRTPWR_c_196_n N_VIRTPWR_c_197_n N_VIRTPWR_c_198_n N_VIRTPWR_c_185_n
+ N_VIRTPWR_c_200_n N_VIRTPWR_c_186_n N_VIRTPWR_c_187_n N_VIRTPWR_c_188_n
+ VIRTPWR N_VIRTPWR_c_189_n PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%VIRTPWR
cc_1 noxref_1 SLEEP 0.058587f $X=-0.19 $Y=-0.002 $X2=8.315 $Y2=0.84
cc_2 noxref_1 N_VPWR_c_92_n 0.618373f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_3 noxref_1 VIRTPWR 0.105802f $X=-0.19 $Y=-0.002 $X2=8.377 $Y2=2.4
cc_4 noxref_1 N_VIRTPWR_c_185_n 0.0836651f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_5 noxref_1 N_VIRTPWR_c_186_n 0.0786895f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_6 noxref_1 N_VIRTPWR_c_187_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_7 noxref_1 N_VIRTPWR_c_188_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_8 noxref_1 N_VIRTPWR_c_189_n 0.0386646f $X=-0.19 $Y=-0.002 $X2=0 $Y2=0
cc_9 VPB N_SLEEP_c_38_n 0.045835f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=1.895
cc_10 VPB N_SLEEP_c_39_n 0.0164013f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.325
cc_11 VPB N_SLEEP_c_40_n 0.045835f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.755
cc_12 VPB N_SLEEP_c_41_n 0.0108874f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=2.325
cc_13 VPB SLEEP 0.0289324f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=0.84
cc_14 VPB N_SLEEP_c_43_n 0.0240095f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=1.985
cc_15 VPB N_SLEEP_c_44_n 0.0240095f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=2.665
cc_16 VPB N_VPWR_c_93_n 0.0994951f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=1.985
cc_17 VPB N_VPWR_c_94_n 0.00214921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_95_n 0.0155703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_96_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_97_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_98_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_99_n 0.00821471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_92_n 0.115514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_24 VPB N_VIRTPWR_c_190_n 0.0130323f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.755
cc_25 VPB N_VIRTPWR_c_191_n 0.0357155f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=2.25
cc_26 VPB N_VIRTPWR_c_192_n 0.15875f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=2.665
cc_27 VPB N_VIRTPWR_c_193_n 0.00789876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VIRTPWR_c_194_n 0.00789876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_VIRTPWR_c_195_n 0.00789876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VIRTPWR_c_196_n 0.00815152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VIRTPWR_c_197_n 0.00214921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VIRTPWR_c_198_n 0.0329627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VIRTPWR_c_185_n 0.0405705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VIRTPWR_c_200_n 0.0130323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_VIRTPWR_c_186_n 0.0404102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 N_SLEEP_c_38_n N_VPWR_c_93_n 0.0112707f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_37 SLEEP N_VPWR_c_93_n 0.0122857f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_38 N_SLEEP_c_39_n N_VPWR_c_94_n 0.0102402f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_39 N_SLEEP_c_40_n N_VPWR_c_94_n 0.010275f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_40 SLEEP N_VPWR_c_94_n 0.0107074f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_41 N_SLEEP_c_44_n N_VPWR_c_94_n 0.00207026f $X=8.42 $Y=2.665 $X2=0 $Y2=0
cc_42 N_SLEEP_c_38_n N_VPWR_c_95_n 0.00410997f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_43 N_SLEEP_c_39_n N_VPWR_c_95_n 0.00343818f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_44 N_SLEEP_c_40_n N_VPWR_c_95_n 0.00303147f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_45 N_SLEEP_c_38_n N_VPWR_c_96_n 0.00101546f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_46 N_SLEEP_c_39_n N_VPWR_c_96_n 0.00101546f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_47 N_SLEEP_c_38_n N_VPWR_c_97_n 0.00101546f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_48 N_SLEEP_c_39_n N_VPWR_c_97_n 0.00101546f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_49 N_SLEEP_c_38_n N_VPWR_c_98_n 0.00101546f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_50 N_SLEEP_c_39_n N_VPWR_c_98_n 0.00101546f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_51 N_SLEEP_c_38_n N_VPWR_c_99_n 0.00320659f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_52 N_SLEEP_c_39_n N_VPWR_c_99_n 0.00320659f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_53 SLEEP N_VPWR_c_99_n 0.0205357f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_54 N_SLEEP_c_38_n N_VPWR_c_92_n 0.00718609f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_55 N_SLEEP_c_39_n N_VPWR_c_92_n 0.00392683f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_56 N_SLEEP_c_40_n N_VPWR_c_92_n 0.00984441f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_57 SLEEP N_VPWR_c_92_n 0.100759f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_58 N_SLEEP_c_43_n N_VPWR_c_92_n 0.00118998f $X=8.42 $Y=1.985 $X2=0 $Y2=0
cc_59 N_SLEEP_c_44_n N_VPWR_c_92_n 0.00118998f $X=8.42 $Y=2.665 $X2=0 $Y2=0
cc_60 N_SLEEP_c_40_n N_VIRTPWR_c_190_n 0.0158929f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_61 N_SLEEP_c_40_n N_VIRTPWR_c_191_n 0.00259154f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_62 N_SLEEP_c_38_n N_VIRTPWR_c_193_n 0.00101539f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_63 N_SLEEP_c_39_n N_VIRTPWR_c_193_n 0.00101539f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_64 N_SLEEP_c_40_n N_VIRTPWR_c_193_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_65 N_SLEEP_c_38_n N_VIRTPWR_c_194_n 0.00101539f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_66 N_SLEEP_c_39_n N_VIRTPWR_c_194_n 0.00101539f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_67 N_SLEEP_c_40_n N_VIRTPWR_c_194_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_68 N_SLEEP_c_38_n N_VIRTPWR_c_195_n 0.00101539f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_69 N_SLEEP_c_39_n N_VIRTPWR_c_195_n 0.00101539f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_70 N_SLEEP_c_40_n N_VIRTPWR_c_195_n 0.00539584f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_71 N_SLEEP_c_38_n N_VIRTPWR_c_196_n 0.00101545f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_72 N_SLEEP_c_39_n N_VIRTPWR_c_196_n 0.00101545f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_73 N_SLEEP_c_40_n N_VIRTPWR_c_196_n 0.00539734f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_74 N_SLEEP_c_38_n N_VIRTPWR_c_197_n 0.0102402f $X=8.17 $Y=1.895 $X2=0 $Y2=0
cc_75 N_SLEEP_c_39_n N_VIRTPWR_c_197_n 0.0102402f $X=8.17 $Y=2.325 $X2=0 $Y2=0
cc_76 SLEEP N_VIRTPWR_c_197_n 0.0107074f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_77 N_SLEEP_c_43_n N_VIRTPWR_c_197_n 0.00207026f $X=8.42 $Y=1.985 $X2=0 $Y2=0
cc_78 N_SLEEP_c_40_n N_VIRTPWR_c_198_n 0.00576677f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_79 SLEEP N_VIRTPWR_c_198_n 0.0165417f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_80 N_SLEEP_c_40_n N_VIRTPWR_c_185_n 0.0037323f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_81 SLEEP N_VIRTPWR_c_185_n 0.0123629f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_82 N_SLEEP_c_40_n N_VIRTPWR_c_186_n 0.00224979f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_83 N_VPWR_c_95_n N_VIRTPWR_M1000_d 3.18208e-19 $X=1.545 $Y=1.68 $X2=-0.19
+ $Y2=-0.002
cc_84 N_VPWR_c_99_n N_VIRTPWR_M1000_d 2.87889e-19 $X=7.775 $Y=1.68 $X2=-0.19
+ $Y2=-0.002
cc_85 N_VPWR_c_94_n N_VIRTPWR_c_190_n 0.262559f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_86 N_VPWR_c_95_n N_VIRTPWR_c_190_n 0.00580238f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_87 N_VPWR_c_92_n N_VIRTPWR_c_190_n 0.00611837f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_88 N_VPWR_c_92_n VIRTPWR 0.224849f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_89 N_VPWR_c_96_n N_VIRTPWR_c_192_n 0.00708574f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_90 N_VPWR_c_97_n N_VIRTPWR_c_192_n 0.00708574f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_91 N_VPWR_c_98_n N_VIRTPWR_c_192_n 0.00708574f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_92 N_VPWR_c_99_n N_VIRTPWR_c_192_n 0.00580238f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_93 N_VPWR_c_92_n N_VIRTPWR_c_192_n 0.0186573f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_94 N_VPWR_M1001_s N_VIRTPWR_c_193_n 2.87738e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_95 N_VPWR_c_93_n N_VIRTPWR_c_193_n 0.0389016f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_96 N_VPWR_c_94_n N_VIRTPWR_c_193_n 0.0346616f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_97 N_VPWR_c_95_n N_VIRTPWR_c_193_n 0.0970367f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_98 N_VPWR_c_96_n N_VIRTPWR_c_193_n 0.0970367f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_99 N_VPWR_c_92_n N_VIRTPWR_c_193_n 0.219944f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_100 N_VPWR_M1001_s N_VIRTPWR_c_194_n 2.87738e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_101 N_VPWR_c_93_n N_VIRTPWR_c_194_n 0.0389016f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_102 N_VPWR_c_94_n N_VIRTPWR_c_194_n 0.0346616f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_103 N_VPWR_c_96_n N_VIRTPWR_c_194_n 0.0970367f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_104 N_VPWR_c_97_n N_VIRTPWR_c_194_n 0.0970367f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_105 N_VPWR_c_92_n N_VIRTPWR_c_194_n 0.219944f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_106 N_VPWR_M1001_s N_VIRTPWR_c_195_n 2.87738e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_107 N_VPWR_c_93_n N_VIRTPWR_c_195_n 0.0389016f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_108 N_VPWR_c_94_n N_VIRTPWR_c_195_n 0.0346616f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_109 N_VPWR_c_97_n N_VIRTPWR_c_195_n 0.0970367f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_110 N_VPWR_c_98_n N_VIRTPWR_c_195_n 0.0970367f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_111 N_VPWR_c_92_n N_VIRTPWR_c_195_n 0.219944f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_112 N_VPWR_M1001_s N_VIRTPWR_c_196_n 2.8786e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_113 N_VPWR_c_93_n N_VIRTPWR_c_196_n 0.0400253f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_114 N_VPWR_c_94_n N_VIRTPWR_c_196_n 0.0356496f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_115 N_VPWR_c_98_n N_VIRTPWR_c_196_n 0.0970546f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_116 N_VPWR_c_99_n N_VIRTPWR_c_196_n 0.0970546f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_117 N_VPWR_c_92_n N_VIRTPWR_c_196_n 0.225341f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_118 N_VPWR_c_93_n N_VIRTPWR_c_197_n 0.251237f $X=7.785 $Y=1.68 $X2=0 $Y2=0
cc_119 N_VPWR_c_94_n N_VIRTPWR_c_197_n 0.251237f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_120 N_VPWR_c_95_n N_VIRTPWR_c_197_n 0.0377876f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_121 N_VPWR_c_96_n N_VIRTPWR_c_197_n 0.0358966f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_122 N_VPWR_c_97_n N_VIRTPWR_c_197_n 0.0358966f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_123 N_VPWR_c_98_n N_VIRTPWR_c_197_n 0.0358966f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_124 N_VPWR_c_99_n N_VIRTPWR_c_197_n 0.0393669f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_125 N_VPWR_c_92_n N_VIRTPWR_c_197_n 0.0173287f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_126 N_VPWR_c_94_n N_VIRTPWR_c_185_n 0.00290716f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_127 N_VPWR_c_99_n N_VIRTPWR_c_185_n 0.026124f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_128 N_VPWR_c_92_n N_VIRTPWR_c_185_n 0.227442f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_129 N_VPWR_c_92_n N_VIRTPWR_c_200_n 0.00787277f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_130 N_VPWR_c_94_n N_VIRTPWR_c_186_n 0.00285709f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_131 N_VPWR_c_95_n N_VIRTPWR_c_186_n 0.026124f $X=1.545 $Y=1.68 $X2=0 $Y2=0
cc_132 N_VPWR_c_92_n N_VIRTPWR_c_186_n 0.212348f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_133 N_VPWR_c_94_n N_VIRTPWR_c_187_n 0.0012824f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_134 N_VPWR_c_96_n N_VIRTPWR_c_187_n 0.0229031f $X=3.09 $Y=1.68 $X2=0 $Y2=0
cc_135 N_VPWR_c_92_n N_VIRTPWR_c_187_n 0.0980574f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_136 N_VPWR_c_94_n N_VIRTPWR_c_188_n 0.0012824f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_137 N_VPWR_c_97_n N_VIRTPWR_c_188_n 0.0229031f $X=4.645 $Y=1.68 $X2=0 $Y2=0
cc_138 N_VPWR_c_92_n N_VIRTPWR_c_188_n 0.0980574f $X=7.775 $Y=1.68 $X2=0 $Y2=0
cc_139 N_VPWR_c_94_n N_VIRTPWR_c_189_n 0.0012824f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_140 N_VPWR_c_98_n N_VIRTPWR_c_189_n 0.0229031f $X=6.2 $Y=1.68 $X2=0 $Y2=0
cc_141 N_VPWR_c_92_n N_VIRTPWR_c_189_n 0.0980574f $X=7.775 $Y=1.68 $X2=0 $Y2=0
