* NGSPICE file created from sky130_fd_sc_lp__or4_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or4_2 A B C D VGND VNB VPB VPWR X
M1000 a_72_367# B VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=9.429e+11p ps=8.24e+06u
M1001 a_335_367# B a_227_367# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.638e+11p ps=1.62e+06u
M1002 VGND C a_72_367# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_72_367# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1004 X a_72_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=8.148e+11p ps=6.8e+06u
M1005 a_227_367# C a_155_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 VGND A a_72_367# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_335_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_155_367# D a_72_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 VPWR a_72_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_72_367# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_72_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

