* File: sky130_fd_sc_lp__nor4bb_lp.spice
* Created: Fri Aug 28 10:59:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4bb_lp.pex.spice"
.subckt sky130_fd_sc_lp__nor4bb_lp  VNB VPB C_N B A D_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D_N	D_N
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1007 A_144_47# N_C_N_M1007_g N_A_27_409#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004.8 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_C_N_M1001_g A_144_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75004.4
+ A=0.063 P=1.14 MULT=1
MM1008 A_302_47# N_A_27_409#_M1008_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75004
+ A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_A_27_409#_M1009_g A_302_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1013 A_460_47# N_A_430_21#_M1013_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_430_21#_M1014_g A_460_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0441 PD=0.73 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1002 A_624_47# N_B_M1002_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0651 PD=0.63 PS=0.73 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75002.6 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g A_624_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003 SB=75002 A=0.063
+ P=1.14 MULT=1
MM1010 A_782_47# N_A_M1010_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0588 PD=0.69 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75003.4 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g A_782_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0567 PD=0.84 PS=0.69 NRD=0 NRS=22.848 M=1 R=2.8 SA=75003.8 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1015 A_980_47# N_D_N_M1015_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=39.996 M=1 R=2.8 SA=75004.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_430_21#_M1017_d N_D_N_M1017_g A_980_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75004.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_C_N_M1005_g N_A_27_409#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1016 N_A_352_409#_M1016_d N_A_27_409#_M1016_g N_A_245_409#_M1016_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1000 N_A_245_409#_M1000_d N_A_430_21#_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1003 A_788_409# N_B_M1003_g N_A_352_409#_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g A_788_409# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.12 PD=1.32 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_A_430_21#_M1006_d N_D_N_M1006_g N_VPWR_M1011_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=7.8603 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.6163 P=16.29
c_101 VPB 0 7.95967e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nor4bb_lp.pxi.spice"
*
.ends
*
*
