* File: sky130_fd_sc_lp__invlp_2.spice
* Created: Wed Sep  2 09:57:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__invlp_2.pex.spice"
.subckt sky130_fd_sc_lp__invlp_2  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_116_55#_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1002 N_A_116_55#_M1001_s N_A_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1007 N_A_116_55#_M1007_d N_A_M1007_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_116_55#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.147 PD=2.25 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_116_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1004 N_A_116_367#_M1000_s N_A_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_A_116_367#_M1005_d N_A_M1005_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_116_367#_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4473 AS=0.1764 PD=3.23 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.3 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__invlp_2.pxi.spice"
*
.ends
*
*
