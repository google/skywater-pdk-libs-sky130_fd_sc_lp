* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_0 A B VGND VNB VPB VPWR X
X0 a_27_481# B a_110_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VGND B a_27_481# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_481# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_110_481# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 X a_27_481# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_317_85# B X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR A a_274_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_274_481# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND A a_317_85# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_27_481# a_274_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
