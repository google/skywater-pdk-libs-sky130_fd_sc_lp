* File: sky130_fd_sc_lp__a41o_0.pex.spice
* Created: Fri Aug 28 10:02:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41O_0%A_80_309# 1 2 8 11 15 17 19 22 23 24 25 28 31
+ 33 34 35 39
c78 34 0 1.8157e-19 $X=0.59 $Y=1.71
c79 24 0 1.36801e-19 $X=1.15 $Y=2.13
r80 36 39 12.4248 $w=3.18e-07 $l=3.45e-07 $layer=LI1_cond $X=1.29 $Y=0.44
+ $X2=1.635 $Y2=0.44
r81 34 42 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.71
+ $X2=0.577 $Y2=1.545
r82 33 35 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=1.71 $X2=0.7
+ $Y2=1.545
r83 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.71 $X2=0.59 $Y2=1.71
r84 30 36 2.18543 $w=2.5e-07 $l=1.6e-07 $layer=LI1_cond $X=1.29 $Y=0.6 $X2=1.29
+ $Y2=0.44
r85 30 31 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.29 $Y=0.6 $X2=1.29
+ $Y2=0.74
r86 26 28 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=1.297 $Y=2.215
+ $X2=1.297 $Y2=2.51
r87 24 26 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.15 $Y=2.13
+ $X2=1.297 $Y2=2.215
r88 24 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.15 $Y=2.13
+ $X2=0.895 $Y2=2.13
r89 22 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.165 $Y=0.825
+ $X2=1.29 $Y2=0.74
r90 22 23 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.165 $Y=0.825
+ $X2=0.895 $Y2=0.825
r91 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.81 $Y=0.91
+ $X2=0.895 $Y2=0.825
r92 20 35 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.81 $Y=0.91
+ $X2=0.81 $Y2=1.545
r93 19 25 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=0.7 $Y=2.045
+ $X2=0.895 $Y2=2.13
r94 18 33 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=0.7 $Y=1.74 $X2=0.7
+ $Y2=1.71
r95 18 19 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=0.7 $Y=1.74 $X2=0.7
+ $Y2=2.045
r96 15 42 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=0.65 $Y=0.445
+ $X2=0.65 $Y2=1.545
r97 11 17 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.475 $Y=2.725
+ $X2=0.475 $Y2=2.215
r98 8 17 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.577 $Y=2.038
+ $X2=0.577 $Y2=2.215
r99 7 34 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=1.722
+ $X2=0.577 $Y2=1.71
r100 7 8 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.577 $Y=1.722
+ $X2=0.577 $Y2=2.038
r101 2 28 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.19
+ $Y=2.365 $X2=1.315 $Y2=2.51
r102 1 39 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.235 $X2=1.635 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%B1 3 6 9 13 14 17 19 20 24
c55 19 0 1.8157e-19 $X=1.2 $Y=1.295
c56 6 0 1.28941e-19 $X=1.25 $Y=2.065
r57 19 20 16.1342 $w=2.98e-07 $l=4.2e-07 $layer=LI1_cond $X=1.215 $Y=1.245
+ $X2=1.215 $Y2=1.665
r58 19 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.245 $X2=1.16 $Y2=1.245
r59 15 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.25 $Y=2.14
+ $X2=1.53 $Y2=2.14
r60 13 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.585
+ $X2=1.16 $Y2=1.245
r61 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.585
+ $X2=1.16 $Y2=1.75
r62 12 24 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.08
+ $X2=1.16 $Y2=1.245
r63 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.53 $Y=2.215
+ $X2=1.53 $Y2=2.14
r64 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.53 $Y=2.215 $X2=1.53
+ $Y2=2.685
r65 6 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.25 $Y=2.065
+ $X2=1.25 $Y2=2.14
r66 6 14 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.25 $Y=2.065
+ $X2=1.25 $Y2=1.75
r67 3 12 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.08 $Y=0.445
+ $X2=1.08 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%A1 5 9 11 12 13 14 15 20
c51 13 0 1.28941e-19 $X=1.68 $Y=0.925
c52 9 0 1.36801e-19 $X=1.96 $Y=2.685
r53 20 22 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=1.32
+ $X2=1.745 $Y2=1.155
r54 14 15 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=1.295
+ $X2=1.717 $Y2=1.665
r55 14 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.32 $X2=1.73 $Y2=1.32
r56 13 14 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.717 $Y=0.925
+ $X2=1.717 $Y2=1.295
r57 11 12 44.1784 $w=3.6e-07 $l=1.5e-07 $layer=POLY_cond $X=1.8 $Y=1.675 $X2=1.8
+ $Y2=1.825
r58 9 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.96 $Y=2.685
+ $X2=1.96 $Y2=1.825
r59 5 22 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.85 $Y=0.445
+ $X2=1.85 $Y2=1.155
r60 1 20 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.745 $Y=1.335
+ $X2=1.745 $Y2=1.32
r61 1 11 54.4984 $w=3.6e-07 $l=3.4e-07 $layer=POLY_cond $X=1.745 $Y=1.335
+ $X2=1.745 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%A2 3 6 9 10 11 12 13 14 15 21
c47 12 0 5.07064e-20 $X=2.16 $Y=0.555
r48 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.3 $Y=0.93
+ $X2=2.3 $Y2=0.93
r49 14 15 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.197 $Y=1.295
+ $X2=2.197 $Y2=1.665
r50 14 22 11.2171 $w=3.73e-07 $l=3.65e-07 $layer=LI1_cond $X=2.197 $Y=1.295
+ $X2=2.197 $Y2=0.93
r51 13 22 0.153659 $w=3.73e-07 $l=5e-09 $layer=LI1_cond $X=2.197 $Y=0.925
+ $X2=2.197 $Y2=0.93
r52 12 13 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.197 $Y=0.555
+ $X2=2.197 $Y2=0.925
r53 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.3 $Y=1.27 $X2=2.3
+ $Y2=0.93
r54 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.27 $X2=2.3
+ $Y2=1.435
r55 9 21 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=0.765 $X2=2.3
+ $Y2=0.93
r56 6 11 640.957 $w=1.5e-07 $l=1.25e-06 $layer=POLY_cond $X=2.39 $Y=2.685
+ $X2=2.39 $Y2=1.435
r57 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.31 $Y=0.445 $X2=2.31
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%A3 3 6 9 11 12 13 14 19
c42 12 0 9.34739e-20 $X=3.12 $Y=0.925
c43 9 0 2.12067e-19 $X=2.82 $Y=2.685
r44 19 21 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.32
+ $X2=2.855 $Y2=1.155
r45 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.87
+ $Y=1.32 $X2=2.87 $Y2=1.32
r46 14 20 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3 $Y=1.665 $X2=3
+ $Y2=1.32
r47 13 20 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3 $Y=1.295 $X2=3
+ $Y2=1.32
r48 12 13 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3 $Y=0.925 $X2=3
+ $Y2=1.295
r49 9 11 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.82 $Y=2.685
+ $X2=2.82 $Y2=1.825
r50 6 11 40.9331 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=2.855 $Y=1.645
+ $X2=2.855 $Y2=1.825
r51 5 19 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=2.855 $Y=1.335
+ $X2=2.855 $Y2=1.32
r52 5 6 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=2.855 $Y=1.335
+ $X2=2.855 $Y2=1.645
r53 3 21 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.75 $Y=0.445
+ $X2=2.75 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%A4 1 3 6 9 13 17 20 21 22 23 28
c39 21 0 4.68024e-20 $X=3.6 $Y=0.925
c40 17 0 9.34739e-20 $X=3.38 $Y=2.14
r41 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.47
+ $Y=1.005 $X2=3.47 $Y2=1.005
r42 22 23 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.665
r43 22 29 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.005
r44 21 29 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=3.57 $Y=0.925 $X2=3.57
+ $Y2=1.005
r45 19 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.47 $Y=1.345
+ $X2=3.47 $Y2=1.005
r46 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.47 $Y=1.345
+ $X2=3.47 $Y2=1.51
r47 15 17 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=3.275 $Y=2.14
+ $X2=3.38 $Y2=2.14
r48 13 28 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.47 $Y=0.915 $X2=3.47
+ $Y2=1.005
r49 10 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.11 $Y=0.84
+ $X2=3.47 $Y2=0.84
r50 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.38 $Y=2.065
+ $X2=3.38 $Y2=2.14
r51 9 20 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.38 $Y=2.065
+ $X2=3.38 $Y2=1.51
r52 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.275 $Y=2.215
+ $X2=3.275 $Y2=2.14
r53 4 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.275 $Y=2.215 $X2=3.275
+ $Y2=2.685
r54 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.11 $Y=0.765
+ $X2=3.11 $Y2=0.84
r55 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.11 $Y=0.765 $X2=3.11
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%X 1 2 7 8 9 10 11 12 13 37 46 49
r18 49 50 1.16452 $w=3.03e-07 $l=2e-08 $layer=LI1_cond $X=0.237 $Y=2.405
+ $X2=0.237 $Y2=2.385
r19 35 37 0.491205 $w=3.03e-07 $l=1.3e-08 $layer=LI1_cond $X=0.237 $Y=2.537
+ $X2=0.237 $Y2=2.55
r20 23 41 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=0.61
+ $X2=0.21 $Y2=0.445
r21 13 37 8.50163 $w=3.03e-07 $l=2.25e-07 $layer=LI1_cond $X=0.237 $Y=2.775
+ $X2=0.237 $Y2=2.55
r22 12 35 3.7785 $w=3.03e-07 $l=1e-07 $layer=LI1_cond $X=0.237 $Y=2.437
+ $X2=0.237 $Y2=2.537
r23 12 49 1.20912 $w=3.03e-07 $l=3.2e-08 $layer=LI1_cond $X=0.237 $Y=2.437
+ $X2=0.237 $Y2=2.405
r24 12 50 1.52122 $w=2.48e-07 $l=3.3e-08 $layer=LI1_cond $X=0.21 $Y=2.352
+ $X2=0.21 $Y2=2.385
r25 11 12 14.613 $w=2.48e-07 $l=3.17e-07 $layer=LI1_cond $X=0.21 $Y=2.035
+ $X2=0.21 $Y2=2.352
r26 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r27 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r28 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=0.925 $X2=0.21
+ $Y2=1.295
r29 7 46 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.24 $Y=0.445
+ $X2=0.435 $Y2=0.445
r30 7 41 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.445 $X2=0.21
+ $Y2=0.445
r31 7 8 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=0.21 $Y=0.625 $X2=0.21
+ $Y2=0.925
r32 7 23 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.21 $Y=0.625
+ $X2=0.21 $Y2=0.61
r33 2 37 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.26 $Y2=2.55
r34 1 46 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.235 $X2=0.435 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%VPWR 1 2 3 12 16 20 23 24 25 27 32 42 43 46
+ 49
r50 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 37 49 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.172 $Y2=3.33
r57 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 36 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 33 46 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.707 $Y2=3.33
r61 33 35 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 32 49 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=2.172 $Y2=3.33
r63 32 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 30 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 27 46 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.707 $Y2=3.33
r67 27 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r68 25 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 25 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 23 39 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=2.64
+ $Y2=3.33
r71 23 24 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=3.045 $Y2=3.33
r72 22 42 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.19 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 22 24 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.19 $Y=3.33
+ $X2=3.045 $Y2=3.33
r74 18 24 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.045 $Y2=3.33
r75 18 20 29.2085 $w=2.88e-07 $l=7.35e-07 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.045 $Y2=2.51
r76 14 49 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.172 $Y=3.245
+ $X2=2.172 $Y2=3.33
r77 14 16 31.964 $w=2.63e-07 $l=7.35e-07 $layer=LI1_cond $X=2.172 $Y=3.245
+ $X2=2.172 $Y2=2.51
r78 10 46 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=3.245
+ $X2=0.707 $Y2=3.33
r79 10 12 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=0.707 $Y=3.245
+ $X2=0.707 $Y2=2.55
r80 3 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.365 $X2=3.035 $Y2=2.51
r81 2 16 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.035
+ $Y=2.365 $X2=2.175 $Y2=2.51
r82 1 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.405 $X2=0.69 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%A_321_473# 1 2 3 12 14 15 18 20 24 26
c45 24 0 1.14558e-19 $X=3.49 $Y=2.51
r46 22 24 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=3.507 $Y=2.175
+ $X2=3.507 $Y2=2.51
r47 21 26 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.73 $Y=2.09
+ $X2=2.602 $Y2=2.09
r48 20 22 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=3.36 $Y=2.09
+ $X2=3.507 $Y2=2.175
r49 20 21 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.36 $Y=2.09
+ $X2=2.73 $Y2=2.09
r50 16 26 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.602 $Y=2.175
+ $X2=2.602 $Y2=2.09
r51 16 18 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=2.602 $Y=2.175
+ $X2=2.602 $Y2=2.51
r52 14 26 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.475 $Y=2.09
+ $X2=2.602 $Y2=2.09
r53 14 15 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.475 $Y=2.09
+ $X2=1.87 $Y2=2.09
r54 10 15 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.742 $Y=2.175
+ $X2=1.87 $Y2=2.09
r55 10 12 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=1.742 $Y=2.175
+ $X2=1.742 $Y2=2.51
r56 3 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.35
+ $Y=2.365 $X2=3.49 $Y2=2.51
r57 2 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=2.365 $X2=2.605 $Y2=2.51
r58 1 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.605
+ $Y=2.365 $X2=1.745 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_0%VGND 1 2 9 13 16 17 19 20 21 34 35
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r52 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r53 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 28 31 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r55 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r57 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 21 32 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r59 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r60 19 31 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.12
+ $Y2=0
r61 19 20 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.332
+ $Y2=0
r62 18 34 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.53 $Y=0 $X2=3.6
+ $Y2=0
r63 18 20 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=3.53 $Y=0 $X2=3.332
+ $Y2=0
r64 16 24 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.72
+ $Y2=0
r65 16 17 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.867
+ $Y2=0
r66 15 28 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.2
+ $Y2=0
r67 15 17 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.867
+ $Y2=0
r68 11 20 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.332 $Y=0.085
+ $X2=3.332 $Y2=0
r69 11 13 10.2115 $w=3.93e-07 $l=3.5e-07 $layer=LI1_cond $X=3.332 $Y=0.085
+ $X2=3.332 $Y2=0.435
r70 7 17 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.867 $Y=0.085
+ $X2=0.867 $Y2=0
r71 7 9 14.462 $w=2.53e-07 $l=3.2e-07 $layer=LI1_cond $X=0.867 $Y=0.085
+ $X2=0.867 $Y2=0.405
r72 2 13 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.235 $X2=3.325 $Y2=0.435
r73 1 9 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.725
+ $Y=0.235 $X2=0.865 $Y2=0.405
.ends

