* File: sky130_fd_sc_lp__mux2i_lp.pxi.spice
* Created: Wed Sep  2 10:01:30 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2I_LP%S N_S_c_70_n N_S_c_85_n N_S_c_86_n N_S_M1001_g
+ N_S_M1010_g N_S_c_72_n N_S_M1003_g N_S_M1011_g N_S_M1000_g N_S_c_75_n
+ N_S_M1004_g N_S_c_76_n N_S_c_77_n N_S_c_93_p N_S_c_167_p N_S_c_78_n N_S_c_79_n
+ N_S_c_80_n N_S_c_81_n S N_S_c_82_n N_S_c_83_n PM_SKY130_FD_SC_LP__MUX2I_LP%S
x_PM_SKY130_FD_SC_LP__MUX2I_LP%A1 N_A1_M1008_g N_A1_M1009_g N_A1_c_185_n
+ N_A1_c_186_n N_A1_c_190_n N_A1_c_191_n A1 N_A1_c_187_n
+ PM_SKY130_FD_SC_LP__MUX2I_LP%A1
x_PM_SKY130_FD_SC_LP__MUX2I_LP%A0 N_A0_M1002_g N_A0_c_256_n N_A0_c_252_n
+ N_A0_M1005_g N_A0_c_254_n A0 A0 N_A0_c_259_n PM_SKY130_FD_SC_LP__MUX2I_LP%A0
x_PM_SKY130_FD_SC_LP__MUX2I_LP%A_365_255# N_A_365_255#_M1004_d
+ N_A_365_255#_M1000_d N_A_365_255#_M1007_g N_A_365_255#_M1006_g
+ N_A_365_255#_c_312_n N_A_365_255#_c_313_n N_A_365_255#_c_314_n
+ N_A_365_255#_c_315_n N_A_365_255#_c_316_n
+ PM_SKY130_FD_SC_LP__MUX2I_LP%A_365_255#
x_PM_SKY130_FD_SC_LP__MUX2I_LP%VPWR N_VPWR_M1010_s N_VPWR_M1007_d N_VPWR_c_376_n
+ N_VPWR_c_377_n N_VPWR_c_378_n VPWR N_VPWR_c_379_n N_VPWR_c_380_n
+ N_VPWR_c_375_n N_VPWR_c_382_n PM_SKY130_FD_SC_LP__MUX2I_LP%VPWR
x_PM_SKY130_FD_SC_LP__MUX2I_LP%Y N_Y_M1008_d N_Y_M1002_d N_Y_c_416_n N_Y_c_414_n
+ N_Y_c_418_n N_Y_c_419_n N_Y_c_420_n N_Y_c_415_n Y Y Y
+ PM_SKY130_FD_SC_LP__MUX2I_LP%Y
x_PM_SKY130_FD_SC_LP__MUX2I_LP%VGND N_VGND_M1001_s N_VGND_M1006_d N_VGND_c_493_n
+ N_VGND_c_494_n N_VGND_c_495_n VGND N_VGND_c_496_n N_VGND_c_497_n
+ N_VGND_c_498_n N_VGND_c_499_n PM_SKY130_FD_SC_LP__MUX2I_LP%VGND
cc_1 VNB N_S_c_70_n 0.0151434f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=2.295
cc_2 VNB N_S_M1001_g 0.0242514f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.455
cc_3 VNB N_S_c_72_n 0.016917f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.775
cc_4 VNB N_S_M1011_g 0.0241877f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.845
cc_5 VNB N_S_M1000_g 0.0296259f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=2.845
cc_6 VNB N_S_c_75_n 0.0196285f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=0.775
cc_7 VNB N_S_c_76_n 0.00513426f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.9
cc_8 VNB N_S_c_77_n 0.00251151f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.815
cc_9 VNB N_S_c_78_n 6.36605e-19 $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=0.775
cc_10 VNB N_S_c_79_n 0.0117247f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.98
cc_11 VNB N_S_c_80_n 0.0927946f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.98
cc_12 VNB N_S_c_81_n 0.00400636f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.94
cc_13 VNB N_S_c_82_n 0.00726219f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=0.94
cc_14 VNB N_S_c_83_n 0.0363352f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=0.94
cc_15 VNB N_A1_M1008_g 0.040253f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.37
cc_16 VNB N_A1_c_185_n 0.00686055f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.845
cc_17 VNB N_A1_c_186_n 0.0104811f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.845
cc_18 VNB N_A1_c_187_n 0.0320835f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=2.845
cc_19 VNB N_A0_c_252_n 0.0328045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A0_M1005_g 0.023251f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.845
cc_21 VNB N_A0_c_254_n 0.011421f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.455
cc_22 VNB N_A_365_255#_M1007_g 0.0028233f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.445
cc_23 VNB N_A_365_255#_M1006_g 0.0411736f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.775
cc_24 VNB N_A_365_255#_c_312_n 0.0211427f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.455
cc_25 VNB N_A_365_255#_c_313_n 0.0280779f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.845
cc_26 VNB N_A_365_255#_c_314_n 0.0021126f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=2.845
cc_27 VNB N_A_365_255#_c_315_n 0.0440736f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=0.455
cc_28 VNB N_A_365_255#_c_316_n 0.0152709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_375_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.86 $Y2=0.455
cc_30 VNB N_Y_c_414_n 0.00648316f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.845
cc_31 VNB N_Y_c_415_n 0.0100974f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=2.845
cc_32 VNB N_VGND_c_493_n 0.0110794f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.455
cc_33 VNB N_VGND_c_494_n 0.0184472f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.445
cc_34 VNB N_VGND_c_495_n 0.00594176f $X=-0.19 $Y=-0.245 $X2=2.47 $Y2=0.775
cc_35 VNB N_VGND_c_496_n 0.0379779f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.845
cc_36 VNB N_VGND_c_497_n 0.0297459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_498_n 0.189531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_499_n 0.00631837f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.34
cc_39 VPB N_S_c_70_n 0.0524361f $X=-0.19 $Y=1.655 $X2=0.18 $Y2=2.295
cc_40 VPB N_S_c_85_n 0.0214047f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.37
cc_41 VPB N_S_c_86_n 0.0154367f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=2.37
cc_42 VPB N_S_M1010_g 0.0272568f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.845
cc_43 VPB N_S_M1011_g 0.0636557f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=2.845
cc_44 VPB N_S_M1000_g 0.0707875f $X=-0.19 $Y=1.655 $X2=2.835 $Y2=2.845
cc_45 VPB N_A1_M1009_g 0.0220145f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.455
cc_46 VPB N_A1_c_185_n 0.007316f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.845
cc_47 VPB N_A1_c_190_n 0.00870127f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=0.455
cc_48 VPB N_A1_c_191_n 0.0294736f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=1.105
cc_49 VPB N_A0_M1002_g 0.0443402f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.37
cc_50 VPB N_A0_c_256_n 0.0358276f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.815
cc_51 VPB N_A0_c_252_n 0.00428883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB A0 0.0150767f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=1.105
cc_53 VPB N_A0_c_259_n 0.0446998f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=0.775
cc_54 VPB N_A_365_255#_M1007_g 0.0636348f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.445
cc_55 VPB N_A_365_255#_c_314_n 0.0619862f $X=-0.19 $Y=1.655 $X2=2.835 $Y2=2.845
cc_56 VPB N_VPWR_c_376_n 0.0130354f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.455
cc_57 VPB N_VPWR_c_377_n 0.024263f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.445
cc_58 VPB N_VPWR_c_378_n 0.00397614f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=0.775
cc_59 VPB N_VPWR_c_379_n 0.042725f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=2.845
cc_60 VPB N_VPWR_c_380_n 0.0276647f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=0.775
cc_61 VPB N_VPWR_c_375_n 0.0736833f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=0.455
cc_62 VPB N_VPWR_c_382_n 0.00540913f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.425
cc_63 VPB N_Y_c_416_n 0.00341055f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.455
cc_64 VPB N_Y_c_414_n 6.49329e-19 $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.845
cc_65 VPB N_Y_c_418_n 0.0137843f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.845
cc_66 VPB N_Y_c_419_n 0.00151901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_Y_c_420_n 0.0050882f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=0.775
cc_68 VPB Y 0.00980503f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=0.775
cc_69 VPB Y 0.00956418f $X=-0.19 $Y=1.655 $X2=2.86 $Y2=0.455
cc_70 N_S_M1001_g N_A1_M1008_g 0.0347137f $X=0.495 $Y=0.455 $X2=0 $Y2=0
cc_71 N_S_c_76_n N_A1_M1008_g 0.0020592f $X=0.615 $Y=0.9 $X2=0 $Y2=0
cc_72 N_S_c_77_n N_A1_M1008_g 0.00217485f $X=0.7 $Y=0.815 $X2=0 $Y2=0
cc_73 N_S_c_93_p N_A1_M1008_g 0.014505f $X=1.72 $Y=0.34 $X2=0 $Y2=0
cc_74 N_S_c_79_n N_A1_M1008_g 8.26796e-19 $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_75 N_S_c_76_n N_A1_c_186_n 0.0157937f $X=0.615 $Y=0.9 $X2=0 $Y2=0
cc_76 N_S_c_79_n N_A1_c_186_n 0.0273718f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_77 N_S_c_80_n N_A1_c_186_n 0.00289566f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_78 N_S_c_79_n N_A1_c_187_n 2.37823e-19 $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_79 N_S_c_80_n N_A1_c_187_n 0.0347137f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_80 N_S_c_70_n N_A0_M1002_g 0.00261396f $X=0.18 $Y=2.295 $X2=0 $Y2=0
cc_81 N_S_c_85_n N_A0_M1002_g 0.0475402f $X=0.475 $Y=2.37 $X2=0 $Y2=0
cc_82 N_S_c_81_n N_A0_c_252_n 4.72313e-19 $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_83 N_S_c_93_p N_A0_M1005_g 0.0124428f $X=1.72 $Y=0.34 $X2=0 $Y2=0
cc_84 N_S_c_78_n N_A0_M1005_g 0.00479882f $X=1.805 $Y=0.775 $X2=0 $Y2=0
cc_85 N_S_c_81_n N_A0_M1005_g 0.00182553f $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_86 N_S_c_70_n A0 0.0350288f $X=0.18 $Y=2.295 $X2=0 $Y2=0
cc_87 N_S_c_85_n A0 0.0101192f $X=0.475 $Y=2.37 $X2=0 $Y2=0
cc_88 N_S_c_79_n A0 0.0198091f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_89 N_S_c_80_n A0 0.00580418f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_90 N_S_c_70_n N_A0_c_259_n 0.0149718f $X=0.18 $Y=2.295 $X2=0 $Y2=0
cc_91 N_S_c_85_n N_A0_c_259_n 0.00500433f $X=0.475 $Y=2.37 $X2=0 $Y2=0
cc_92 N_S_c_80_n N_A0_c_259_n 0.00217096f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_93 N_S_M1011_g N_A_365_255#_M1007_g 0.0344377f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_94 N_S_c_72_n N_A_365_255#_M1006_g 0.0237259f $X=2.47 $Y=0.775 $X2=0 $Y2=0
cc_95 N_S_M1011_g N_A_365_255#_M1006_g 0.00636088f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_96 N_S_c_93_p N_A_365_255#_M1006_g 0.00380777f $X=1.72 $Y=0.34 $X2=0 $Y2=0
cc_97 N_S_c_78_n N_A_365_255#_M1006_g 0.00727133f $X=1.805 $Y=0.775 $X2=0 $Y2=0
cc_98 N_S_c_81_n N_A_365_255#_M1006_g 0.00346617f $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_99 N_S_c_82_n N_A_365_255#_M1006_g 0.013059f $X=2.56 $Y=0.94 $X2=0 $Y2=0
cc_100 N_S_M1011_g N_A_365_255#_c_312_n 0.0202501f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_101 N_S_M1000_g N_A_365_255#_c_312_n 0.0186639f $X=2.835 $Y=2.845 $X2=0 $Y2=0
cc_102 N_S_c_81_n N_A_365_255#_c_312_n 0.00534641f $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_103 N_S_c_82_n N_A_365_255#_c_312_n 0.0659323f $X=2.56 $Y=0.94 $X2=0 $Y2=0
cc_104 N_S_c_83_n N_A_365_255#_c_312_n 8.1708e-19 $X=2.835 $Y=0.94 $X2=0 $Y2=0
cc_105 N_S_M1011_g N_A_365_255#_c_313_n 0.0176381f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_106 N_S_c_81_n N_A_365_255#_c_313_n 9.53394e-19 $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_107 N_S_c_82_n N_A_365_255#_c_313_n 0.00330343f $X=2.56 $Y=0.94 $X2=0 $Y2=0
cc_108 N_S_M1011_g N_A_365_255#_c_314_n 0.00495933f $X=2.475 $Y=2.845 $X2=0
+ $Y2=0
cc_109 N_S_M1000_g N_A_365_255#_c_314_n 0.0483356f $X=2.835 $Y=2.845 $X2=0 $Y2=0
cc_110 N_S_c_72_n N_A_365_255#_c_315_n 0.00184301f $X=2.47 $Y=0.775 $X2=0 $Y2=0
cc_111 N_S_c_75_n N_A_365_255#_c_315_n 0.0117654f $X=2.86 $Y=0.775 $X2=0 $Y2=0
cc_112 N_S_c_82_n N_A_365_255#_c_315_n 0.0251958f $X=2.56 $Y=0.94 $X2=0 $Y2=0
cc_113 N_S_c_83_n N_A_365_255#_c_315_n 0.0192896f $X=2.835 $Y=0.94 $X2=0 $Y2=0
cc_114 N_S_M1000_g N_A_365_255#_c_316_n 0.0088642f $X=2.835 $Y=2.845 $X2=0 $Y2=0
cc_115 N_S_c_86_n N_VPWR_c_377_n 0.00797826f $X=0.255 $Y=2.37 $X2=0 $Y2=0
cc_116 N_S_M1010_g N_VPWR_c_377_n 0.0145258f $X=0.55 $Y=2.845 $X2=0 $Y2=0
cc_117 N_S_M1011_g N_VPWR_c_378_n 0.0103146f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_118 N_S_M1000_g N_VPWR_c_378_n 0.00168354f $X=2.835 $Y=2.845 $X2=0 $Y2=0
cc_119 N_S_M1010_g N_VPWR_c_379_n 0.00452967f $X=0.55 $Y=2.845 $X2=0 $Y2=0
cc_120 N_S_M1011_g N_VPWR_c_380_n 0.00452967f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_121 N_S_M1000_g N_VPWR_c_380_n 0.00511358f $X=2.835 $Y=2.845 $X2=0 $Y2=0
cc_122 N_S_c_86_n N_VPWR_c_375_n 0.00164531f $X=0.255 $Y=2.37 $X2=0 $Y2=0
cc_123 N_S_M1010_g N_VPWR_c_375_n 0.00809218f $X=0.55 $Y=2.845 $X2=0 $Y2=0
cc_124 N_S_M1011_g N_VPWR_c_375_n 0.00799963f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_125 N_S_M1000_g N_VPWR_c_375_n 0.0102504f $X=2.835 $Y=2.845 $X2=0 $Y2=0
cc_126 N_S_c_93_p N_Y_M1008_d 0.0102408f $X=1.72 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_127 N_S_c_76_n N_Y_c_414_n 0.00209313f $X=0.615 $Y=0.9 $X2=0 $Y2=0
cc_128 N_S_c_81_n N_Y_c_414_n 0.0144878f $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_129 N_S_M1011_g N_Y_c_418_n 0.0025991f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_130 N_S_c_81_n N_Y_c_418_n 0.0036171f $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_131 N_S_M1010_g N_Y_c_420_n 0.00130204f $X=0.55 $Y=2.845 $X2=0 $Y2=0
cc_132 N_S_c_76_n N_Y_c_415_n 0.00729349f $X=0.615 $Y=0.9 $X2=0 $Y2=0
cc_133 N_S_c_77_n N_Y_c_415_n 0.011114f $X=0.7 $Y=0.815 $X2=0 $Y2=0
cc_134 N_S_c_93_p N_Y_c_415_n 0.0313826f $X=1.72 $Y=0.34 $X2=0 $Y2=0
cc_135 N_S_c_78_n N_Y_c_415_n 0.0138308f $X=1.805 $Y=0.775 $X2=0 $Y2=0
cc_136 N_S_c_81_n N_Y_c_415_n 0.0129541f $X=1.89 $Y=0.94 $X2=0 $Y2=0
cc_137 N_S_M1011_g Y 0.00594528f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_138 N_S_M1011_g Y 0.0044109f $X=2.475 $Y=2.845 $X2=0 $Y2=0
cc_139 N_S_M1001_g N_VGND_c_494_n 0.0105681f $X=0.495 $Y=0.455 $X2=0 $Y2=0
cc_140 N_S_c_76_n N_VGND_c_494_n 6.36887e-19 $X=0.615 $Y=0.9 $X2=0 $Y2=0
cc_141 N_S_c_79_n N_VGND_c_494_n 0.0245598f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_142 N_S_c_80_n N_VGND_c_494_n 0.00220605f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_143 N_S_c_72_n N_VGND_c_495_n 0.00327461f $X=2.47 $Y=0.775 $X2=0 $Y2=0
cc_144 N_S_c_82_n N_VGND_c_495_n 0.0250467f $X=2.56 $Y=0.94 $X2=0 $Y2=0
cc_145 N_S_M1001_g N_VGND_c_496_n 0.00477554f $X=0.495 $Y=0.455 $X2=0 $Y2=0
cc_146 N_S_c_93_p N_VGND_c_496_n 0.0630672f $X=1.72 $Y=0.34 $X2=0 $Y2=0
cc_147 N_S_c_167_p N_VGND_c_496_n 0.0104206f $X=0.785 $Y=0.34 $X2=0 $Y2=0
cc_148 N_S_c_72_n N_VGND_c_497_n 0.00575161f $X=2.47 $Y=0.775 $X2=0 $Y2=0
cc_149 N_S_c_75_n N_VGND_c_497_n 0.00539298f $X=2.86 $Y=0.775 $X2=0 $Y2=0
cc_150 N_S_c_83_n N_VGND_c_497_n 0.00110773f $X=2.835 $Y=0.94 $X2=0 $Y2=0
cc_151 N_S_M1001_g N_VGND_c_498_n 0.00444075f $X=0.495 $Y=0.455 $X2=0 $Y2=0
cc_152 N_S_c_72_n N_VGND_c_498_n 0.00613773f $X=2.47 $Y=0.775 $X2=0 $Y2=0
cc_153 N_S_c_75_n N_VGND_c_498_n 0.0108283f $X=2.86 $Y=0.775 $X2=0 $Y2=0
cc_154 N_S_c_76_n N_VGND_c_498_n 0.00514203f $X=0.615 $Y=0.9 $X2=0 $Y2=0
cc_155 N_S_c_93_p N_VGND_c_498_n 0.0402527f $X=1.72 $Y=0.34 $X2=0 $Y2=0
cc_156 N_S_c_167_p N_VGND_c_498_n 0.00660921f $X=0.785 $Y=0.34 $X2=0 $Y2=0
cc_157 N_S_c_79_n N_VGND_c_498_n 0.00148812f $X=0.27 $Y=0.98 $X2=0 $Y2=0
cc_158 N_S_c_82_n N_VGND_c_498_n 0.0181149f $X=2.56 $Y=0.94 $X2=0 $Y2=0
cc_159 N_S_c_83_n N_VGND_c_498_n 0.00150372f $X=2.835 $Y=0.94 $X2=0 $Y2=0
cc_160 N_S_c_77_n A_114_49# 2.57545e-19 $X=0.7 $Y=0.815 $X2=-0.19 $Y2=-0.245
cc_161 N_S_c_167_p A_114_49# 0.00126025f $X=0.785 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_162 N_S_c_93_p A_324_49# 0.00280851f $X=1.72 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_163 N_S_c_78_n A_324_49# 0.00246143f $X=1.805 $Y=0.775 $X2=-0.19 $Y2=-0.245
cc_164 N_A1_M1009_g N_A0_M1002_g 0.0173024f $X=1.37 $Y=2.845 $X2=0 $Y2=0
cc_165 N_A1_c_190_n N_A0_M1002_g 0.00933517f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_166 N_A1_c_191_n N_A0_M1002_g 0.0162383f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_167 N_A1_c_185_n N_A0_c_256_n 0.012158f $X=1.12 $Y=2.115 $X2=0 $Y2=0
cc_168 N_A1_c_190_n N_A0_c_256_n 0.00347007f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_169 N_A1_c_191_n N_A0_c_256_n 0.0183346f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_170 N_A1_c_185_n N_A0_c_252_n 0.00146594f $X=1.12 $Y=2.115 $X2=0 $Y2=0
cc_171 N_A1_c_186_n N_A0_c_252_n 0.00115023f $X=1.035 $Y=1.32 $X2=0 $Y2=0
cc_172 N_A1_c_187_n N_A0_c_252_n 0.0139557f $X=0.975 $Y=1.32 $X2=0 $Y2=0
cc_173 N_A1_M1008_g N_A0_M1005_g 0.0156112f $X=0.885 $Y=0.455 $X2=0 $Y2=0
cc_174 N_A1_M1008_g N_A0_c_254_n 0.0053675f $X=0.885 $Y=0.455 $X2=0 $Y2=0
cc_175 N_A1_c_185_n A0 0.030485f $X=1.12 $Y=2.115 $X2=0 $Y2=0
cc_176 N_A1_c_186_n A0 0.0159713f $X=1.035 $Y=1.32 $X2=0 $Y2=0
cc_177 N_A1_c_190_n A0 0.00289313f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_178 N_A1_c_187_n A0 2.34807e-19 $X=0.975 $Y=1.32 $X2=0 $Y2=0
cc_179 N_A1_c_185_n N_A0_c_259_n 0.0065622f $X=1.12 $Y=2.115 $X2=0 $Y2=0
cc_180 N_A1_c_186_n N_A0_c_259_n 0.00593421f $X=1.035 $Y=1.32 $X2=0 $Y2=0
cc_181 N_A1_c_187_n N_A0_c_259_n 0.0195695f $X=0.975 $Y=1.32 $X2=0 $Y2=0
cc_182 N_A1_M1009_g N_A_365_255#_M1007_g 0.0221212f $X=1.37 $Y=2.845 $X2=0 $Y2=0
cc_183 N_A1_c_185_n N_A_365_255#_M1007_g 0.00105788f $X=1.12 $Y=2.115 $X2=0
+ $Y2=0
cc_184 N_A1_c_190_n N_A_365_255#_M1007_g 3.67398e-19 $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_185 N_A1_c_191_n N_A_365_255#_M1007_g 0.0180844f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_186 N_A1_M1009_g N_VPWR_c_379_n 0.00373561f $X=1.37 $Y=2.845 $X2=0 $Y2=0
cc_187 N_A1_M1009_g N_VPWR_c_375_n 0.00550909f $X=1.37 $Y=2.845 $X2=0 $Y2=0
cc_188 N_A1_M1009_g N_Y_c_416_n 0.0091177f $X=1.37 $Y=2.845 $X2=0 $Y2=0
cc_189 N_A1_c_190_n N_Y_c_416_n 0.0194485f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_190 N_A1_c_191_n N_Y_c_416_n 0.00313888f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_191 N_A1_M1008_g N_Y_c_414_n 0.0032847f $X=0.885 $Y=0.455 $X2=0 $Y2=0
cc_192 N_A1_c_185_n N_Y_c_414_n 0.0209448f $X=1.12 $Y=2.115 $X2=0 $Y2=0
cc_193 N_A1_c_186_n N_Y_c_414_n 0.0270169f $X=1.035 $Y=1.32 $X2=0 $Y2=0
cc_194 N_A1_c_187_n N_Y_c_414_n 8.98809e-19 $X=0.975 $Y=1.32 $X2=0 $Y2=0
cc_195 N_A1_c_190_n N_Y_c_418_n 0.00259285f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_196 N_A1_c_185_n N_Y_c_419_n 0.0132329f $X=1.12 $Y=2.115 $X2=0 $Y2=0
cc_197 N_A1_c_190_n N_Y_c_419_n 0.01429f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_198 N_A1_c_191_n N_Y_c_419_n 0.00115173f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_199 N_A1_M1009_g N_Y_c_420_n 0.00795856f $X=1.37 $Y=2.845 $X2=0 $Y2=0
cc_200 N_A1_c_190_n N_Y_c_420_n 0.0239582f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_201 N_A1_c_191_n N_Y_c_420_n 9.19985e-19 $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_202 N_A1_M1008_g N_Y_c_415_n 0.00374021f $X=0.885 $Y=0.455 $X2=0 $Y2=0
cc_203 N_A1_c_186_n N_Y_c_415_n 0.0106652f $X=1.035 $Y=1.32 $X2=0 $Y2=0
cc_204 N_A1_c_187_n N_Y_c_415_n 6.33248e-19 $X=0.975 $Y=1.32 $X2=0 $Y2=0
cc_205 N_A1_c_185_n Y 0.00617375f $X=1.12 $Y=2.115 $X2=0 $Y2=0
cc_206 N_A1_c_190_n Y 0.0204015f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_207 N_A1_c_191_n Y 8.715e-19 $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_208 N_A1_M1009_g Y 0.0038579f $X=1.37 $Y=2.845 $X2=0 $Y2=0
cc_209 N_A1_c_190_n Y 0.0076503f $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_210 N_A1_c_191_n Y 3.25253e-19 $X=1.42 $Y=2.28 $X2=0 $Y2=0
cc_211 N_A1_M1008_g N_VGND_c_494_n 0.00130662f $X=0.885 $Y=0.455 $X2=0 $Y2=0
cc_212 N_A1_M1008_g N_VGND_c_496_n 0.00351226f $X=0.885 $Y=0.455 $X2=0 $Y2=0
cc_213 N_A1_M1008_g N_VGND_c_498_n 0.00571852f $X=0.885 $Y=0.455 $X2=0 $Y2=0
cc_214 N_A0_c_256_n N_A_365_255#_M1007_g 0.0157237f $X=1.435 $Y=1.8 $X2=0 $Y2=0
cc_215 N_A0_c_252_n N_A_365_255#_M1006_g 0.0106044f $X=1.51 $Y=1.725 $X2=0 $Y2=0
cc_216 N_A0_M1005_g N_A_365_255#_M1006_g 0.0476373f $X=1.545 $Y=0.455 $X2=0
+ $Y2=0
cc_217 N_A0_c_252_n N_A_365_255#_c_312_n 0.00106799f $X=1.51 $Y=1.725 $X2=0
+ $Y2=0
cc_218 N_A0_c_252_n N_A_365_255#_c_313_n 0.0157237f $X=1.51 $Y=1.725 $X2=0 $Y2=0
cc_219 N_A0_M1002_g N_VPWR_c_377_n 0.00216401f $X=0.94 $Y=2.845 $X2=0 $Y2=0
cc_220 A0 N_VPWR_c_377_n 0.0141451f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_221 N_A0_M1002_g N_VPWR_c_379_n 0.00511358f $X=0.94 $Y=2.845 $X2=0 $Y2=0
cc_222 N_A0_M1002_g N_VPWR_c_375_n 0.00961121f $X=0.94 $Y=2.845 $X2=0 $Y2=0
cc_223 N_A0_c_256_n N_Y_c_414_n 0.00334491f $X=1.435 $Y=1.8 $X2=0 $Y2=0
cc_224 N_A0_c_252_n N_Y_c_414_n 0.0203664f $X=1.51 $Y=1.725 $X2=0 $Y2=0
cc_225 N_A0_c_254_n N_Y_c_414_n 0.00317313f $X=1.527 $Y=1.035 $X2=0 $Y2=0
cc_226 N_A0_c_256_n N_Y_c_418_n 0.00299665f $X=1.435 $Y=1.8 $X2=0 $Y2=0
cc_227 N_A0_c_256_n N_Y_c_419_n 0.00377948f $X=1.435 $Y=1.8 $X2=0 $Y2=0
cc_228 N_A0_M1002_g N_Y_c_420_n 0.00981185f $X=0.94 $Y=2.845 $X2=0 $Y2=0
cc_229 N_A0_M1005_g N_Y_c_415_n 0.00979674f $X=1.545 $Y=0.455 $X2=0 $Y2=0
cc_230 N_A0_c_254_n N_Y_c_415_n 0.00232562f $X=1.527 $Y=1.035 $X2=0 $Y2=0
cc_231 N_A0_M1005_g N_VGND_c_496_n 0.00351226f $X=1.545 $Y=0.455 $X2=0 $Y2=0
cc_232 N_A0_M1005_g N_VGND_c_498_n 0.00571852f $X=1.545 $Y=0.455 $X2=0 $Y2=0
cc_233 N_A_365_255#_M1007_g N_VPWR_c_378_n 0.0100365f $X=1.9 $Y=2.845 $X2=0
+ $Y2=0
cc_234 N_A_365_255#_c_314_n N_VPWR_c_378_n 0.00975716f $X=3.05 $Y=2.845 $X2=0
+ $Y2=0
cc_235 N_A_365_255#_M1007_g N_VPWR_c_379_n 0.00387722f $X=1.9 $Y=2.845 $X2=0
+ $Y2=0
cc_236 N_A_365_255#_c_314_n N_VPWR_c_380_n 0.0252211f $X=3.05 $Y=2.845 $X2=0
+ $Y2=0
cc_237 N_A_365_255#_M1007_g N_VPWR_c_375_n 0.00595485f $X=1.9 $Y=2.845 $X2=0
+ $Y2=0
cc_238 N_A_365_255#_c_314_n N_VPWR_c_375_n 0.013614f $X=3.05 $Y=2.845 $X2=0
+ $Y2=0
cc_239 N_A_365_255#_M1006_g N_Y_c_414_n 0.00116459f $X=1.935 $Y=0.455 $X2=0
+ $Y2=0
cc_240 N_A_365_255#_c_312_n N_Y_c_414_n 0.0169814f $X=2.885 $Y=1.44 $X2=0 $Y2=0
cc_241 N_A_365_255#_c_313_n N_Y_c_414_n 0.00142409f $X=1.99 $Y=1.44 $X2=0 $Y2=0
cc_242 N_A_365_255#_M1007_g N_Y_c_418_n 0.00940122f $X=1.9 $Y=2.845 $X2=0 $Y2=0
cc_243 N_A_365_255#_c_312_n N_Y_c_418_n 0.0377691f $X=2.885 $Y=1.44 $X2=0 $Y2=0
cc_244 N_A_365_255#_c_313_n N_Y_c_418_n 0.00433126f $X=1.99 $Y=1.44 $X2=0 $Y2=0
cc_245 N_A_365_255#_c_314_n N_Y_c_418_n 0.00544132f $X=3.05 $Y=2.845 $X2=0 $Y2=0
cc_246 N_A_365_255#_M1007_g N_Y_c_420_n 0.00143436f $X=1.9 $Y=2.845 $X2=0 $Y2=0
cc_247 N_A_365_255#_M1006_g N_Y_c_415_n 2.91717e-19 $X=1.935 $Y=0.455 $X2=0
+ $Y2=0
cc_248 N_A_365_255#_M1007_g Y 0.0148213f $X=1.9 $Y=2.845 $X2=0 $Y2=0
cc_249 N_A_365_255#_c_314_n Y 0.0127601f $X=3.05 $Y=2.845 $X2=0 $Y2=0
cc_250 N_A_365_255#_M1007_g Y 0.0190835f $X=1.9 $Y=2.845 $X2=0 $Y2=0
cc_251 N_A_365_255#_c_314_n Y 0.00812838f $X=3.05 $Y=2.845 $X2=0 $Y2=0
cc_252 N_A_365_255#_M1006_g N_VGND_c_495_n 0.00501109f $X=1.935 $Y=0.455 $X2=0
+ $Y2=0
cc_253 N_A_365_255#_M1006_g N_VGND_c_496_n 0.00530333f $X=1.935 $Y=0.455 $X2=0
+ $Y2=0
cc_254 N_A_365_255#_c_315_n N_VGND_c_497_n 0.0210519f $X=3.075 $Y=0.47 $X2=0
+ $Y2=0
cc_255 N_A_365_255#_M1004_d N_VGND_c_498_n 0.00229188f $X=2.935 $Y=0.245 $X2=0
+ $Y2=0
cc_256 N_A_365_255#_M1006_g N_VGND_c_498_n 0.00611948f $X=1.935 $Y=0.455 $X2=0
+ $Y2=0
cc_257 N_A_365_255#_c_315_n N_VGND_c_498_n 0.0126421f $X=3.075 $Y=0.47 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_379_n N_Y_c_416_n 0.00870178f $X=2.095 $Y=3.33 $X2=0 $Y2=0
cc_259 N_VPWR_c_375_n N_Y_c_416_n 0.0126955f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_c_377_n N_Y_c_420_n 0.0145731f $X=0.335 $Y=2.845 $X2=0 $Y2=0
cc_261 N_VPWR_c_379_n N_Y_c_420_n 0.0226753f $X=2.095 $Y=3.33 $X2=0 $Y2=0
cc_262 N_VPWR_c_375_n N_Y_c_420_n 0.0124056f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_263 N_VPWR_c_378_n Y 0.0157208f $X=2.26 $Y=2.89 $X2=0 $Y2=0
cc_264 N_VPWR_c_379_n Y 0.00606951f $X=2.095 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_c_375_n Y 0.0104393f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_266 N_Y_c_416_n A_289_527# 0.00408261f $X=1.755 $Y=2.7 $X2=-0.19 $Y2=-0.245
cc_267 Y A_289_527# 2.11515e-19 $X=2.075 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_268 N_Y_M1008_d N_VGND_c_498_n 0.00410159f $X=0.96 $Y=0.245 $X2=0 $Y2=0
cc_269 N_VGND_c_498_n A_114_49# 0.00221166f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_270 N_VGND_c_498_n A_324_49# 0.00193007f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_271 N_VGND_c_498_n A_509_49# 0.00503583f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
