* NGSPICE file created from sky130_fd_sc_lp__a211oi_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a211oi_0 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_148_47# A2 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.289e+11p ps=2.77e+06u
M1001 VGND B1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.717e+11p ps=3.45e+06u
M1002 a_312_483# B1 a_57_483# VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=3.488e+11p ps=3.65e+06u
M1003 VPWR A2 a_57_483# VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1004 Y C1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_57_483# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 a_312_483# VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1007 Y A1 a_148_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

