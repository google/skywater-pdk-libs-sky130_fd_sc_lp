* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_116_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_33_47# B a_116_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR B a_33_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_302_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_302_47# a_33_47# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND B a_302_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_385_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_33_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR A a_385_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 Y a_33_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
