* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 VGND a_27_79# a_196_79# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_1272_128# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_308_463# a_196_79# a_637_191# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_637_191# a_811_341# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 VPWR RESET_B a_1444_320# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND RESET_B a_427_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_861_191# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_811_341# a_27_79# a_1272_128# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_784_191# a_811_341# a_861_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_637_191# a_811_341# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 Q_N a_1272_128# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_811_341# a_196_79# a_1272_128# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_2028_367# a_1272_128# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_308_463# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_637_191# a_27_79# a_793_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_793_463# a_811_341# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VPWR RESET_B a_637_191# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_27_79# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1424_128# a_1444_320# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_79# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_2028_367# a_1272_128# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1582_128# a_1272_128# a_1444_320# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR a_27_79# a_196_79# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_1272_128# a_27_79# a_1424_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR D a_308_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VGND a_2028_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_1272_128# a_196_79# a_1402_496# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 a_1402_496# a_1444_320# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 Q a_2028_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 VGND RESET_B a_1582_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VPWR a_2028_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 VGND a_1272_128# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_308_463# a_27_79# a_637_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 Q_N a_1272_128# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_637_191# a_196_79# a_784_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1444_320# a_1272_128# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X36 a_427_191# D a_308_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 Q a_2028_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
