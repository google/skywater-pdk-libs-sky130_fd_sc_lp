* File: sky130_fd_sc_lp__dlclkp_1.spice
* Created: Fri Aug 28 10:24:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlclkp_1.pex.spice"
.subckt sky130_fd_sc_lp__dlclkp_1  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_80_269#_M1008_g N_A_27_367#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.22485 AS=0.2226 PD=1.84 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1002 A_279_81# N_GATE_M1002_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.112425 PD=0.63 PS=0.92 NRD=14.28 NRS=55.704 M=1 R=2.8
+ SA=75000.9 SB=75002 A=0.063 P=1.14 MULT=1
MM1016 N_A_80_269#_M1016_d N_A_321_55#_M1016_g A_279_81# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1010 A_437_81# N_A_315_382#_M1010_g N_A_80_269#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_27_367#_M1004_g A_437_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0672 PD=0.81 PS=0.74 NRD=24.276 NRS=30 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_A_315_382#_M1012_d N_A_321_55#_M1012_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=7.14 M=1 R=2.8 SA=75002.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_CLK_M1013_g N_A_321_55#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1766 AS=0.1197 PD=1.425 PS=1.41 NRD=104.412 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1007 A_1002_79# N_CLK_M1007_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1766 PD=0.63 PS=1.425 NRD=14.28 NRS=34.284 M=1 R=2.8 SA=75000.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_1046_367#_M1005_d N_A_27_367#_M1005_g A_1002_79# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_GCLK_M1014_d N_A_1046_367#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1019 N_VPWR_M1019_d N_A_80_269#_M1019_g N_A_27_367#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.393385 AS=0.3339 PD=2.55316 PS=3.05 NRD=2.3443 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1018 A_273_480# N_GATE_M1018_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.199815 PD=0.85 PS=1.29684 NRD=15.3857 NRS=114.654 M=1 R=4.26667
+ SA=75001 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1000 N_A_80_269#_M1000_d N_A_315_382#_M1000_g A_273_480# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=12.2928 NRS=15.3857 M=1
+ R=4.26667 SA=75001.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1009 A_453_480# N_A_321_55#_M1009_g N_A_80_269#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0880019 PD=0.63 PS=0.816226 NRD=23.443 NRS=32.8202 M=1
+ R=2.8 SA=75001.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_27_367#_M1001_g A_453_480# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.188346 AS=0.0441 PD=1.23623 PS=0.63 NRD=56.2829 NRS=23.443 M=1 R=2.8
+ SA=75002.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_315_382#_M1003_d N_A_321_55#_M1003_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2752 AS=0.287004 PD=2.14 PS=1.88377 NRD=50.7866 NRS=121.096
+ M=1 R=4.26667 SA=75001.3 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_CLK_M1011_g N_A_321_55#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2365 AS=0.2464 PD=1.74 PS=2.05 NRD=96.8058 NRS=30.7714 M=1
+ R=4.26667 SA=75000.3 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1006 N_A_1046_367#_M1006_d N_CLK_M1006_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2365 PD=0.92 PS=1.74 NRD=0 NRS=96.8058 M=1 R=4.26667
+ SA=75000.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1017 N_VPWR_M1017_d N_A_27_367#_M1017_g N_A_1046_367#_M1006_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.169465 AS=0.0896 PD=1.19242 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001.3 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1015 N_GCLK_M1015_d N_A_1046_367#_M1015_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.333635 PD=3.05 PS=2.34758 NRD=0 NRS=17.9664 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.2415 P=17.93
c_148 VPB 0 7.97162e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlclkp_1.pxi.spice"
*
.ends
*
*
