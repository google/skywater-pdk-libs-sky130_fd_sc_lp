* File: sky130_fd_sc_lp__nand2_lp2.pex.spice
* Created: Fri Aug 28 10:47:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_LP2%B 3 7 9 10 14 15
r29 14 17 65.7961 $w=5.35e-07 $l=5.05e-07 $layer=POLY_cond $X=0.487 $Y=1.275
+ $X2=0.487 $Y2=1.78
r30 14 16 47.5561 $w=5.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.487 $Y=1.275
+ $X2=0.487 $Y2=1.11
r31 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.275 $X2=0.385 $Y2=1.275
r32 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r33 9 15 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.275
r34 7 16 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.68 $Y=0.495
+ $X2=0.68 $Y2=1.11
r35 3 17 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.63 $Y=2.545
+ $X2=0.63 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP2%A 3 5 7 11 12 15 16
r36 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.015 $X2=1.16 $Y2=1.015
r37 12 16 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.16 $Y=1.295
+ $X2=1.16 $Y2=1.015
r38 11 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.355
+ $X2=1.16 $Y2=1.015
r39 10 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=0.85
+ $X2=1.16 $Y2=1.015
r40 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.52
+ $X2=1.16 $Y2=1.355
r41 5 7 254.665 $w=2.5e-07 $l=1.025e-06 $layer=POLY_cond $X=1.16 $Y=1.52
+ $X2=1.16 $Y2=2.545
r42 3 10 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=1.07 $Y=0.495
+ $X2=1.07 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP2%VPWR 1 2 7 9 15 20 21 22 29 30
r23 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 27 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r27 24 33 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.265 $Y2=3.33
r28 24 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.53 $Y=3.33 $X2=1.2
+ $Y2=3.33
r29 22 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r30 22 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 20 26 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.26 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=3.33
+ $X2=1.425 $Y2=3.33
r33 19 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=3.33 $X2=1.68
+ $Y2=3.33
r34 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.59 $Y=3.33
+ $X2=1.425 $Y2=3.33
r35 15 18 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.425 $Y=2.215
+ $X2=1.425 $Y2=2.9
r36 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.425 $Y=3.245
+ $X2=1.425 $Y2=3.33
r37 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.425 $Y=3.245
+ $X2=1.425 $Y2=2.9
r38 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.365 $Y=2.19
+ $X2=0.365 $Y2=2.9
r39 7 33 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.365 $Y=3.245
+ $X2=0.265 $Y2=3.33
r40 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.365 $Y=3.245
+ $X2=0.365 $Y2=2.9
r41 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.285
+ $Y=2.045 $X2=1.425 $Y2=2.9
r42 2 15 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=1.285
+ $Y=2.045 $X2=1.425 $Y2=2.215
r43 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=2.045 $X2=0.365 $Y2=2.9
r44 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=2.045 $X2=0.365 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP2%Y 1 2 9 13 14 16 17 18
r33 18 27 1.14734 $w=3.19e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=0.467 $X2=1.71
+ $Y2=0.467
r34 18 24 15.1066 $w=3.19e-07 $l=3.95e-07 $layer=LI1_cond $X=1.68 $Y=0.467
+ $X2=1.285 $Y2=0.467
r35 17 24 3.25078 $w=3.19e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.467
+ $X2=1.285 $Y2=0.467
r36 15 27 4.42298 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=1.71 $Y=0.67
+ $X2=1.71 $Y2=0.467
r37 15 16 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=1.71 $Y=0.67
+ $X2=1.71 $Y2=1.7
r38 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.625 $Y=1.785
+ $X2=1.71 $Y2=1.7
r39 13 14 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.625 $Y=1.785
+ $X2=1.06 $Y2=1.785
r40 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.895 $Y=2.19
+ $X2=0.895 $Y2=2.9
r41 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.895 $Y=1.87
+ $X2=1.06 $Y2=1.785
r42 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.895 $Y=1.87
+ $X2=0.895 $Y2=2.19
r43 2 11 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=2.045 $X2=0.895 $Y2=2.9
r44 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=2.045 $X2=0.895 $Y2=2.19
r45 1 24 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.285 $X2=1.285 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP2%VGND 1 6 9 10 11 20 21
r17 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r18 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r19 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r20 15 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r21 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r22 11 21 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r23 11 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r24 9 14 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.24 $Y2=0
r25 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.465
+ $Y2=0
r26 8 17 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.72
+ $Y2=0
r27 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.465
+ $Y2=0
r28 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.465 $Y=0.085
+ $X2=0.465 $Y2=0
r29 4 6 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.465 $Y=0.085
+ $X2=0.465 $Y2=0.495
r30 1 6 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.32
+ $Y=0.285 $X2=0.465 $Y2=0.495
.ends

