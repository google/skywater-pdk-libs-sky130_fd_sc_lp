* File: sky130_fd_sc_lp__dlygate4s50_1.spice
* Created: Fri Aug 28 10:30:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlygate4s50_1.pex.spice"
.subckt sky130_fd_sc_lp__dlygate4s50_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_52#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_A_288_52#_M1005_d N_A_27_52#_M1005_g N_VGND_M1003_d VNB NSHORT L=0.5
+ W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=15.708 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1004 N_VGND_M1004_d N_A_288_52#_M1004_g N_A_405_136#_M1004_s VNB NSHORT L=0.5
+ W=0.42 AD=0.0847 AS=0.1113 PD=0.786667 PS=1.37 NRD=18.564 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1000 N_X_M1000_d N_A_405_136#_M1000_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1694 PD=2.21 PS=1.57333 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_27_52#_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=21.0987 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_288_52#_M1006_d N_A_27_52#_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.5
+ W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=30.4759 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1007 N_VPWR_M1007_d N_A_288_52#_M1007_g N_A_405_136#_M1007_s VPB PHIGHVT L=0.5
+ W=0.42 AD=0.09135 AS=0.1113 PD=0.8 PS=1.37 NRD=30.4759 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_X_M1001_d N_A_405_136#_M1001_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.27405 PD=3.05 PS=2.4 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_33 VNB 0 1.65637e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dlygate4s50_1.pxi.spice"
*
.ends
*
*
