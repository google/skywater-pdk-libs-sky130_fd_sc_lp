* File: sky130_fd_sc_lp__a21boi_lp.pex.spice
* Created: Fri Aug 28 09:50:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%A2 3 7 9 10 18
r28 16 18 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.595 $Y=0.975
+ $X2=0.785 $Y2=0.975
r29 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=0.975 $X2=0.595 $Y2=0.975
r30 13 16 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.555 $Y=0.975
+ $X2=0.595 $Y2=0.975
r31 10 17 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.72 $Y=0.975
+ $X2=0.595 $Y2=0.975
r32 9 17 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=0.975
+ $X2=0.595 $Y2=0.975
r33 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.785 $Y=0.81
+ $X2=0.785 $Y2=0.975
r34 5 7 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.785 $Y=0.81
+ $X2=0.785 $Y2=0.445
r35 1 13 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.14
+ $X2=0.555 $Y2=0.975
r36 1 3 349.077 $w=2.5e-07 $l=1.405e-06 $layer=POLY_cond $X=0.555 $Y=1.14
+ $X2=0.555 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%A1 3 7 9 10 11 16
c38 3 0 1.0508e-19 $X=1.085 $Y=2.545
r39 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.625
+ $X2=1.085 $Y2=1.46
r40 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.625 $X2=1.085 $Y2=1.625
r41 11 17 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.625
+ $X2=1.085 $Y2=1.625
r42 10 17 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.72 $Y=1.625
+ $X2=1.085 $Y2=1.625
r43 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.625
+ $X2=0.72 $Y2=1.625
r44 7 18 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=1.175 $Y=0.445
+ $X2=1.175 $Y2=1.46
r45 1 16 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.79
+ $X2=1.085 $Y2=1.625
r46 1 3 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.085 $Y=1.79
+ $X2=1.085 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%A_298_318# 1 2 9 13 15 16 19 24 27 30 31
+ 33 34 37 42 44 47
r81 44 46 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.065 $Y=0.455
+ $X2=3.065 $Y2=0.645
r82 42 47 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.145 $Y=1.675
+ $X2=3.065 $Y2=1.76
r83 42 46 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.145 $Y=1.675
+ $X2=3.145 $Y2=0.645
r84 37 39 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.065 $Y=2.19
+ $X2=3.065 $Y2=2.9
r85 35 47 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=1.845
+ $X2=3.065 $Y2=1.76
r86 35 37 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.065 $Y=1.845
+ $X2=3.065 $Y2=2.19
r87 33 47 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=1.76
+ $X2=3.065 $Y2=1.76
r88 33 34 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.9 $Y=1.76
+ $X2=2.215 $Y2=1.76
r89 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.01
+ $Y=1.235 $X2=2.01 $Y2=1.235
r90 28 34 26.4971 $w=8.2e-08 $l=2.23495e-07 $layer=LI1_cond $X=2.03 $Y=1.675
+ $X2=2.215 $Y2=1.76
r91 28 30 13.7047 $w=3.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.03 $Y=1.675
+ $X2=2.03 $Y2=1.235
r92 26 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.01 $Y=1.22
+ $X2=2.01 $Y2=1.235
r93 26 27 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=2.01 $Y=1.22
+ $X2=2.01 $Y2=1.145
r94 24 31 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.01 $Y=1.59
+ $X2=2.01 $Y2=1.235
r95 17 27 13.5877 $w=2.4e-07 $l=9.48683e-08 $layer=POLY_cond $X=1.965 $Y=1.07
+ $X2=2.01 $Y2=1.145
r96 17 19 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.965 $Y=1.07
+ $X2=1.965 $Y2=0.445
r97 15 27 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.145
+ $X2=2.01 $Y2=1.145
r98 15 16 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.145
+ $X2=1.68 $Y2=1.145
r99 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.605 $Y=1.07
+ $X2=1.68 $Y2=1.145
r100 11 13 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.605 $Y=1.07
+ $X2=1.605 $Y2=0.445
r101 7 24 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.615 $Y=1.665
+ $X2=2.01 $Y2=1.665
r102 7 9 200.005 $w=2.5e-07 $l=8.05e-07 $layer=POLY_cond $X=1.615 $Y=1.74
+ $X2=1.615 $Y2=2.545
r103 2 39 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=2.045 $X2=3.065 $Y2=2.9
r104 2 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=2.045 $X2=3.065 $Y2=2.19
r105 1 44 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.925
+ $Y=0.235 $X2=3.065 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%B1_N 3 7 9 13 15 16 19 20
r41 19 21 82.4947 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=2.67 $Y=0.99
+ $X2=2.67 $Y2=1.495
r42 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.69
+ $Y=0.99 $X2=2.69 $Y2=0.99
r43 16 20 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.69 $Y=1.295
+ $X2=2.69 $Y2=0.99
r44 15 21 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.75 $Y=1.735
+ $X2=2.75 $Y2=1.495
r45 11 19 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.85 $Y=0.825
+ $X2=2.67 $Y2=0.99
r46 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.85 $Y=0.825
+ $X2=2.85 $Y2=0.445
r47 7 15 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.8 $Y=1.86 $X2=2.8
+ $Y2=1.735
r48 7 9 170.191 $w=2.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.8 $Y=1.86 $X2=2.8
+ $Y2=2.545
r49 1 19 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.49 $Y=0.825
+ $X2=2.67 $Y2=0.99
r50 1 3 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.49 $Y=0.825 $X2=2.49
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%A_29_409# 1 2 9 11 16 20
c25 9 0 1.0508e-19 $X=0.29 $Y=2.9
r26 16 18 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.29 $Y=2.19
+ $X2=0.29 $Y2=2.415
r27 12 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=2.415
+ $X2=0.29 $Y2=2.415
r28 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=2.415
+ $X2=1.35 $Y2=2.415
r29 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.185 $Y=2.415
+ $X2=0.455 $Y2=2.415
r30 7 18 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=2.5 $X2=0.29
+ $Y2=2.415
r31 7 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.29 $Y=2.5 $X2=0.29
+ $Y2=2.9
r32 2 20 300 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_PDIFF $count=2 $X=1.21
+ $Y=2.045 $X2=1.35 $Y2=2.495
r33 1 16 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.045 $X2=0.29 $Y2=2.19
r34 1 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.045 $X2=0.29 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%VPWR 1 2 11 15 20 21 22 32 33 36
r38 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r44 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r46 24 26 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 22 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 20 29 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.535 $Y2=3.33
r51 19 32 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.7 $Y=3.33 $X2=3.12
+ $Y2=3.33
r52 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=3.33
+ $X2=2.535 $Y2=3.33
r53 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.535 $Y=2.19
+ $X2=2.535 $Y2=2.9
r54 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=3.245
+ $X2=2.535 $Y2=3.33
r55 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.535 $Y=3.245
+ $X2=2.535 $Y2=2.9
r56 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245 $X2=0.82
+ $Y2=3.33
r57 9 11 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.87
r58 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.045 $X2=2.535 $Y2=2.9
r59 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.045 $X2=2.535 $Y2=2.19
r60 1 11 600 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=2.045 $X2=0.82 $Y2=2.87
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%Y 1 2 8 11 18 20
r41 20 22 6.25641 $w=1.95e-07 $l=1e-07 $layer=LI1_cond $X=1.68 $Y=2.035 $X2=1.58
+ $Y2=2.035
r42 16 18 5.34059 $w=4.08e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=0.47
+ $X2=1.58 $Y2=0.47
r43 11 13 23.3781 $w=3.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.87 $Y=2.19
+ $X2=1.87 $Y2=2.9
r44 9 20 11.8872 $w=1.95e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=2.035
+ $X2=1.68 $Y2=2.035
r45 9 11 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=1.87 $Y=2.15 $X2=1.87
+ $Y2=2.19
r46 8 22 1.54022 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.58 $Y=1.92 $X2=1.58
+ $Y2=2.035
r47 7 18 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.58 $Y=0.675
+ $X2=1.58 $Y2=0.47
r48 7 8 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=1.58 $Y=0.675
+ $X2=1.58 $Y2=1.92
r49 2 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=2.045 $X2=1.88 $Y2=2.9
r50 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=2.045 $X2=1.88 $Y2=2.19
r51 1 16 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.25
+ $Y=0.235 $X2=1.39 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r46 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.18
+ $Y2=0
r48 27 29 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=3.12
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.57
+ $Y2=0
r50 23 25 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.735 $Y=0 $X2=1.68
+ $Y2=0
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=2.18
+ $Y2=0
r52 22 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=1.68
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.405 $Y=0 $X2=0.57
+ $Y2=0
r56 17 19 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.405 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 15 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r59 15 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r61 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0.445
r62 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.57 $Y=0.085 $X2=0.57
+ $Y2=0
r63 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.57 $Y=0.085 $X2=0.57
+ $Y2=0.42
r64 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.18 $Y2=0.445
r65 1 9 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.425
+ $Y=0.235 $X2=0.57 $Y2=0.42
.ends

