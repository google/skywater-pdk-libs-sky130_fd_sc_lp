* File: sky130_fd_sc_lp__dlrtn_4.spice
* Created: Fri Aug 28 10:26:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtn_4.pex.spice"
.subckt sky130_fd_sc_lp__dlrtn_4  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_D_M1016_g N_A_27_468#_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_250_70#_M1001_d N_GATE_N_M1001_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_250_70#_M1017_g N_A_357_365#_M1017_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1003 A_567_125# N_A_27_468#_M1003_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=25.704 M=1 R=2.8 SA=75000.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1024 N_A_639_125#_M1024_d N_A_250_70#_M1024_g A_567_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 A_725_125# N_A_357_365#_M1000_g N_A_639_125#_M1024_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_789_99#_M1004_g A_725_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1018 A_1009_47# N_A_639_125#_M1018_g N_A_789_99#_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_1009_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1785 AS=0.0882 PD=1.265 PS=1.05 NRD=9.276 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1011 N_Q_M1011_d N_A_789_99#_M1011_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1785 PD=1.12 PS=1.265 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1012 N_Q_M1011_d N_A_789_99#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1021 N_Q_M1021_d N_A_789_99#_M1021_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1023 N_Q_M1021_d N_A_789_99#_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 N_VPWR_M1022_d N_D_M1022_g N_A_27_468#_M1022_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.176 AS=0.1696 PD=1.19 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_250_70#_M1005_d N_GATE_N_M1005_g N_VPWR_M1022_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.176 PD=1.81 PS=1.19 NRD=0 NRS=83.0946 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A_250_70#_M1002_g N_A_357_365#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1248 AS=0.3329 PD=1.03 PS=2.82 NRD=16.9223 NRS=143.18 M=1
+ R=4.26667 SA=75000.3 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1010 A_567_447# N_A_27_468#_M1010_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1248 PD=0.85 PS=1.03 NRD=15.3857 NRS=16.9223 M=1 R=4.26667
+ SA=75000.8 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1013 N_A_639_125#_M1013_d N_A_357_365#_M1013_g A_567_447# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.138023 AS=0.0672 PD=1.24981 PS=0.85 NRD=13.0808 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1020 A_748_447# N_A_250_70#_M1020_g N_A_639_125#_M1013_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0905774 PD=0.63 PS=0.820189 NRD=23.443 NRS=35.1645 M=1
+ R=2.8 SA=75001.7 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_789_99#_M1008_g A_748_447# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.139125 AS=0.0441 PD=1.0275 PS=0.63 NRD=129.567 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1019 N_A_789_99#_M1019_d N_A_639_125#_M1019_g N_VPWR_M1008_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.417375 PD=1.54 PS=3.0825 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_RESET_B_M1006_g N_A_789_99#_M1019_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.21735 AS=0.1764 PD=1.605 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4
+ SA=75001.6 SB=75002 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1006_d N_A_789_99#_M1007_g N_Q_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.21735 AS=0.1827 PD=1.605 PS=1.55 NRD=5.4569 NRS=1.5563 M=1 R=8.4
+ SA=75002.1 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_789_99#_M1014_g N_Q_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1827 PD=1.54 PS=1.55 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1014_d N_A_789_99#_M1015_g N_Q_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_A_789_99#_M1025_g N_Q_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=15.0403 P=19.87
c_91 VNB 0 4.62649e-19 $X=0 $Y=0
c_160 VPB 0 8.72356e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlrtn_4.pxi.spice"
*
.ends
*
*
