* File: sky130_fd_sc_lp__srsdfstp_1.pxi.spice
* Created: Wed Sep  2 10:39:22 2020
* 
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%SCD N_SCD_M1001_g N_SCD_M1000_g N_SCD_c_360_n
+ N_SCD_c_365_n SCD SCD N_SCD_c_362_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%SCD
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%D N_D_M1016_g N_D_M1012_g D N_D_c_395_n
+ N_D_c_396_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%D
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_339_93# N_A_339_93#_M1029_s
+ N_A_339_93#_M1036_s N_A_339_93#_M1023_g N_A_339_93#_M1048_g
+ N_A_339_93#_c_434_n N_A_339_93#_c_435_n N_A_339_93#_c_436_n
+ N_A_339_93#_c_437_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_339_93#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%SCE N_SCE_c_483_n N_SCE_M1013_g N_SCE_M1042_g
+ N_SCE_c_485_n N_SCE_c_486_n N_SCE_M1036_g N_SCE_M1029_g N_SCE_c_489_n
+ N_SCE_c_495_n SCE N_SCE_c_491_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%SCE
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_689_139# N_A_689_139#_M1028_d
+ N_A_689_139#_M1010_d N_A_689_139#_c_567_n N_A_689_139#_c_589_n
+ N_A_689_139#_c_590_n N_A_689_139#_c_568_n N_A_689_139#_M1031_g
+ N_A_689_139#_M1005_g N_A_689_139#_M1025_g N_A_689_139#_M1017_g
+ N_A_689_139#_M1021_g N_A_689_139#_c_571_n N_A_689_139#_c_572_n
+ N_A_689_139#_c_573_n N_A_689_139#_c_574_n N_A_689_139#_c_575_n
+ N_A_689_139#_c_576_n N_A_689_139#_c_647_p N_A_689_139#_c_701_p
+ N_A_689_139#_c_596_n N_A_689_139#_c_577_n N_A_689_139#_c_578_n
+ N_A_689_139#_c_597_n N_A_689_139#_c_598_n N_A_689_139#_c_599_n
+ N_A_689_139#_c_724_p N_A_689_139#_c_600_n N_A_689_139#_c_579_n
+ N_A_689_139#_c_601_n N_A_689_139#_c_602_n N_A_689_139#_c_603_n
+ N_A_689_139#_c_580_n N_A_689_139#_c_581_n N_A_689_139#_c_582_n
+ N_A_689_139#_c_583_n N_A_689_139#_c_584_n N_A_689_139#_c_585_n
+ N_A_689_139#_c_609_n N_A_689_139#_c_725_p N_A_689_139#_c_610_n
+ N_A_689_139#_c_586_n N_A_689_139#_c_587_n N_A_689_139#_c_588_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_689_139#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_659_113# N_A_659_113#_M1015_s
+ N_A_659_113#_M1039_d N_A_659_113#_c_896_n N_A_659_113#_M1028_g
+ N_A_659_113#_c_897_n N_A_659_113#_M1010_g N_A_659_113#_c_898_n
+ N_A_659_113#_c_899_n N_A_659_113#_c_900_n N_A_659_113#_M1047_g
+ N_A_659_113#_c_901_n N_A_659_113#_M1034_g N_A_659_113#_c_930_n
+ N_A_659_113#_M1030_g N_A_659_113#_c_931_n N_A_659_113#_c_932_n
+ N_A_659_113#_c_933_n N_A_659_113#_M1037_g N_A_659_113#_c_934_n
+ N_A_659_113#_M1050_g N_A_659_113#_c_936_n N_A_659_113#_c_904_n
+ N_A_659_113#_c_937_n N_A_659_113#_c_938_n N_A_659_113#_c_905_n
+ N_A_659_113#_c_906_n N_A_659_113#_c_907_n N_A_659_113#_c_908_n
+ N_A_659_113#_c_909_n N_A_659_113#_c_910_n N_A_659_113#_c_911_n
+ N_A_659_113#_c_912_n N_A_659_113#_c_913_n N_A_659_113#_c_914_n
+ N_A_659_113#_c_915_n N_A_659_113#_c_916_n N_A_659_113#_c_917_n
+ N_A_659_113#_c_918_n N_A_659_113#_c_939_n N_A_659_113#_c_940_n
+ N_A_659_113#_c_919_n N_A_659_113#_c_920_n N_A_659_113#_c_921_n
+ N_A_659_113#_c_1112_p N_A_659_113#_c_922_n N_A_659_113#_c_923_n
+ N_A_659_113#_c_924_n N_A_659_113#_c_925_n N_A_659_113#_c_926_n
+ N_A_659_113#_c_927_n N_A_659_113#_c_944_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_659_113#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1068_21# N_A_1068_21#_M1038_s
+ N_A_1068_21#_M1009_d N_A_1068_21#_c_1248_n N_A_1068_21#_M1002_g
+ N_A_1068_21#_c_1249_n N_A_1068_21#_c_1250_n N_A_1068_21#_M1035_g
+ N_A_1068_21#_c_1251_n N_A_1068_21#_c_1252_n N_A_1068_21#_c_1256_n
+ N_A_1068_21#_c_1253_n N_A_1068_21#_c_1257_n N_A_1068_21#_c_1258_n
+ N_A_1068_21#_c_1259_n N_A_1068_21#_c_1254_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1068_21#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_887_139# N_A_887_139#_M1047_d
+ N_A_887_139#_M1005_d N_A_887_139#_M1009_g N_A_887_139#_M1038_g
+ N_A_887_139#_M1040_g N_A_887_139#_M1032_g N_A_887_139#_c_1345_n
+ N_A_887_139#_c_1352_n N_A_887_139#_c_1353_n N_A_887_139#_c_1354_n
+ N_A_887_139#_c_1355_n N_A_887_139#_c_1356_n N_A_887_139#_c_1357_n
+ N_A_887_139#_c_1346_n N_A_887_139#_c_1347_n N_A_887_139#_c_1359_n
+ N_A_887_139#_c_1360_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_887_139#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1972_99# N_A_1972_99#_M1041_d
+ N_A_1972_99#_M1018_s N_A_1972_99#_M1046_g N_A_1972_99#_c_1474_n
+ N_A_1972_99#_c_1475_n N_A_1972_99#_M1006_g N_A_1972_99#_c_1477_n
+ N_A_1972_99#_c_1486_n N_A_1972_99#_M1011_g N_A_1972_99#_c_1478_n
+ N_A_1972_99#_c_1479_n N_A_1972_99#_c_1488_n N_A_1972_99#_c_1489_n
+ N_A_1972_99#_c_1531_n N_A_1972_99#_c_1480_n N_A_1972_99#_c_1481_n
+ N_A_1972_99#_c_1491_n N_A_1972_99#_c_1492_n N_A_1972_99#_c_1493_n
+ N_A_1972_99#_c_1482_n N_A_1972_99#_c_1483_n N_A_1972_99#_c_1484_n
+ N_A_1972_99#_c_1485_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1972_99#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_2216_99# N_A_2216_99#_M1022_d
+ N_A_2216_99#_M1045_d N_A_2216_99#_c_1616_n N_A_2216_99#_M1044_g
+ N_A_2216_99#_c_1617_n N_A_2216_99#_c_1618_n N_A_2216_99#_M1024_g
+ N_A_2216_99#_c_1620_n N_A_2216_99#_c_1621_n N_A_2216_99#_c_1622_n
+ N_A_2216_99#_c_1623_n N_A_2216_99#_c_1624_n N_A_2216_99#_c_1625_n
+ N_A_2216_99#_c_1626_n N_A_2216_99#_c_1627_n N_A_2216_99#_c_1628_n
+ N_A_2216_99#_c_1629_n N_A_2216_99#_c_1630_n N_A_2216_99#_c_1631_n
+ N_A_2216_99#_c_1632_n N_A_2216_99#_c_1633_n N_A_2216_99#_c_1634_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_2216_99#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1728_125# N_A_1728_125#_M1017_d
+ N_A_1728_125#_M1037_d N_A_1728_125#_M1043_d N_A_1728_125#_c_1791_n
+ N_A_1728_125#_c_1792_n N_A_1728_125#_c_1793_n N_A_1728_125#_M1051_g
+ N_A_1728_125#_c_1795_n N_A_1728_125#_M1018_g N_A_1728_125#_M1041_g
+ N_A_1728_125#_c_1784_n N_A_1728_125#_c_1785_n N_A_1728_125#_c_1786_n
+ N_A_1728_125#_c_1797_n N_A_1728_125#_c_1798_n N_A_1728_125#_M1019_g
+ N_A_1728_125#_M1007_g N_A_1728_125#_c_1799_n N_A_1728_125#_c_1800_n
+ N_A_1728_125#_c_1823_n N_A_1728_125#_c_1825_n N_A_1728_125#_c_1801_n
+ N_A_1728_125#_c_1830_n N_A_1728_125#_c_1802_n N_A_1728_125#_c_1803_n
+ N_A_1728_125#_c_1833_n N_A_1728_125#_c_1788_n N_A_1728_125#_c_1805_n
+ N_A_1728_125#_c_1844_n N_A_1728_125#_c_1847_n N_A_1728_125#_c_1849_n
+ N_A_1728_125#_c_1789_n N_A_1728_125#_c_1790_n N_A_1728_125#_c_1808_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1728_125#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%SET_B N_SET_B_M1003_g N_SET_B_M1027_g
+ N_SET_B_c_2001_n N_SET_B_c_2002_n N_SET_B_M1008_g N_SET_B_c_2004_n
+ N_SET_B_M1043_g N_SET_B_c_2005_n N_SET_B_c_2006_n N_SET_B_c_2007_n
+ N_SET_B_c_2008_n N_SET_B_c_2009_n SET_B N_SET_B_c_2011_n N_SET_B_c_2012_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%SET_B
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%CLK N_CLK_M1015_g N_CLK_M1039_g CLK CLK CLK
+ N_CLK_c_2123_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%CLK
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%SLEEP_B N_SLEEP_B_M1014_g N_SLEEP_B_M1026_g
+ N_SLEEP_B_M1049_g N_SLEEP_B_c_2171_n N_SLEEP_B_M1045_g N_SLEEP_B_M1020_g
+ N_SLEEP_B_M1022_g N_SLEEP_B_c_2167_n SLEEP_B SLEEP_B N_SLEEP_B_c_2168_n
+ N_SLEEP_B_c_2169_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%SLEEP_B
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_3466_403# N_A_3466_403#_M1007_s
+ N_A_3466_403#_M1019_s N_A_3466_403#_M1004_g N_A_3466_403#_M1033_g
+ N_A_3466_403#_c_2247_n N_A_3466_403#_c_2248_n N_A_3466_403#_c_2239_n
+ N_A_3466_403#_c_2240_n N_A_3466_403#_c_2241_n N_A_3466_403#_c_2242_n
+ N_A_3466_403#_c_2243_n N_A_3466_403#_c_2244_n N_A_3466_403#_c_2245_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_3466_403#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_27_481# N_A_27_481#_M1000_s
+ N_A_27_481#_M1048_d N_A_27_481#_c_2300_n N_A_27_481#_c_2301_n
+ N_A_27_481#_c_2302_n N_A_27_481#_c_2303_n N_A_27_481#_c_2304_n
+ N_A_27_481#_c_2305_n N_A_27_481#_c_2306_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_27_481#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%VPWR N_VPWR_M1000_d N_VPWR_M1036_d
+ N_VPWR_M1035_d N_VPWR_M1027_d N_VPWR_M1019_d N_VPWR_c_2355_n N_VPWR_c_2356_n
+ N_VPWR_c_2357_n N_VPWR_c_2358_n N_VPWR_c_2359_n N_VPWR_c_2360_n
+ N_VPWR_c_2361_n VPWR N_VPWR_c_2362_n N_VPWR_c_2363_n N_VPWR_c_2364_n
+ N_VPWR_c_2365_n N_VPWR_c_2366_n N_VPWR_c_2354_n N_VPWR_c_2368_n
+ N_VPWR_c_2369_n N_VPWR_c_2370_n N_VPWR_c_2371_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_189_119# N_A_189_119#_M1013_d
+ N_A_189_119#_M1047_s N_A_189_119#_M1012_d N_A_189_119#_M1005_s
+ N_A_189_119#_c_2519_n N_A_189_119#_c_2526_n N_A_189_119#_c_2527_n
+ N_A_189_119#_c_2528_n N_A_189_119#_c_2529_n N_A_189_119#_c_2520_n
+ N_A_189_119#_c_2521_n N_A_189_119#_c_2522_n N_A_189_119#_c_2523_n
+ N_A_189_119#_c_2524_n N_A_189_119#_c_2531_n N_A_189_119#_c_2525_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_189_119#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1541_125# N_A_1541_125#_M1040_d
+ N_A_1541_125#_M1032_d N_A_1541_125#_c_2636_n N_A_1541_125#_c_2637_n
+ N_A_1541_125#_c_2653_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_1541_125#
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%KAPWR N_KAPWR_M1018_d N_KAPWR_M1011_d
+ N_KAPWR_M1026_d N_KAPWR_c_2675_n KAPWR N_KAPWR_c_2676_n N_KAPWR_c_2677_n
+ N_KAPWR_c_2678_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%KAPWR
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%Q N_Q_M1033_d N_Q_M1004_d Q Q Q Q Q Q Q
+ N_Q_c_2818_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%Q
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%VGND N_VGND_M1001_s N_VGND_M1023_d
+ N_VGND_M1029_d N_VGND_M1002_d N_VGND_M1003_d N_VGND_M1008_d N_VGND_M1051_s
+ N_VGND_M1049_d N_VGND_M1007_d N_VGND_c_2832_n N_VGND_c_2833_n N_VGND_c_2834_n
+ N_VGND_c_2835_n N_VGND_c_2836_n N_VGND_c_2837_n N_VGND_c_2838_n
+ N_VGND_c_2839_n N_VGND_c_2840_n N_VGND_c_2841_n N_VGND_c_2842_n
+ N_VGND_c_2843_n N_VGND_c_2844_n N_VGND_c_2845_n N_VGND_c_2846_n
+ N_VGND_c_2847_n N_VGND_c_2848_n VGND N_VGND_c_2849_n N_VGND_c_2850_n
+ N_VGND_c_2851_n N_VGND_c_2852_n N_VGND_c_2853_n N_VGND_c_2854_n
+ N_VGND_c_2855_n N_VGND_c_2856_n N_VGND_c_2857_n N_VGND_c_2858_n
+ N_VGND_c_2859_n PM_SKY130_FD_SC_LP__SRSDFSTP_1%VGND
x_PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_2074_125# N_A_2074_125#_M1006_d
+ N_A_2074_125#_M1044_d N_A_2074_125#_c_3022_n N_A_2074_125#_c_3023_n
+ N_A_2074_125#_c_3024_n N_A_2074_125#_c_3025_n
+ PM_SKY130_FD_SC_LP__SRSDFSTP_1%A_2074_125#
cc_1 VNB N_SCD_M1001_g 0.0272437f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.805
cc_2 VNB N_SCD_c_360_n 0.0209451f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.71
cc_3 VNB SCD 0.027856f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_SCD_c_362_n 0.0168098f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_5 VNB N_D_M1016_g 0.0389902f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.805
cc_6 VNB N_D_c_395_n 0.012667f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.875
cc_7 VNB N_D_c_396_n 0.00134235f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_339_93#_M1023_g 0.0272224f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_9 VNB N_A_339_93#_c_434_n 0.00636453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_339_93#_c_435_n 0.0133184f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_11 VNB N_A_339_93#_c_436_n 0.0450718f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_12 VNB N_A_339_93#_c_437_n 0.00825785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_c_483_n 0.0171211f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.805
cc_14 VNB N_SCE_M1013_g 0.0308131f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.725
cc_15 VNB N_SCE_c_485_n 0.15084f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.71
cc_16 VNB N_SCE_c_486_n 0.0125534f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.875
cc_17 VNB N_SCE_M1036_g 6.12425e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCE_M1029_g 0.0376248f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_19 VNB N_SCE_c_489_n 0.0111059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB SCE 0.010715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SCE_c_491_n 0.0387189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_689_139#_c_567_n 0.063754f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.725
cc_23 VNB N_A_689_139#_c_568_n 0.0161165f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.71
cc_24 VNB N_A_689_139#_M1025_g 0.0167653f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_25 VNB N_A_689_139#_M1017_g 0.0206233f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_26 VNB N_A_689_139#_c_571_n 0.0105547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_689_139#_c_572_n 0.0147759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_689_139#_c_573_n 0.0120431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_689_139#_c_574_n 0.00166173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_689_139#_c_575_n 0.0308794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_689_139#_c_576_n 2.76804e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_689_139#_c_577_n 0.00521532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_689_139#_c_578_n 3.26207e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_689_139#_c_579_n 0.0110071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_689_139#_c_580_n 0.00548668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_689_139#_c_581_n 0.00173205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_689_139#_c_582_n 8.74691e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_689_139#_c_583_n 0.0379658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_689_139#_c_584_n 0.00146458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_689_139#_c_585_n 0.003693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_689_139#_c_586_n 0.00377139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_689_139#_c_587_n 0.0105936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_689_139#_c_588_n 0.0609618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_659_113#_c_896_n 0.0201325f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.725
cc_45 VNB N_A_659_113#_c_897_n 0.011605f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.205
cc_46 VNB N_A_659_113#_c_898_n 0.0449863f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_47 VNB N_A_659_113#_c_899_n 0.0152826f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_48 VNB N_A_659_113#_c_900_n 0.0184144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_659_113#_c_901_n 0.0733355f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_50 VNB N_A_659_113#_M1034_g 0.0124437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_659_113#_M1050_g 0.0491575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_659_113#_c_904_n 0.00597897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_659_113#_c_905_n 0.00360532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_659_113#_c_906_n 0.0293673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_659_113#_c_907_n 0.00301202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_659_113#_c_908_n 0.00246568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_659_113#_c_909_n 0.00582445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_659_113#_c_910_n 0.0135878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_659_113#_c_911_n 0.00353283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_659_113#_c_912_n 0.00427867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_659_113#_c_913_n 0.00709532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_659_113#_c_914_n 0.00255969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_659_113#_c_915_n 0.00376091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_659_113#_c_916_n 0.0629219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_659_113#_c_917_n 0.00157725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_659_113#_c_918_n 0.00762158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_659_113#_c_919_n 0.0210419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_659_113#_c_920_n 0.00380715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_659_113#_c_921_n 0.00275359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_659_113#_c_922_n 0.010159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_659_113#_c_923_n 0.0226804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_659_113#_c_924_n 0.00822805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_659_113#_c_925_n 0.0084953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_659_113#_c_926_n 8.84711e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_659_113#_c_927_n 0.00456904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1068_21#_c_1248_n 0.0200642f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.725
cc_77 VNB N_A_1068_21#_c_1249_n 0.0314128f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.205
cc_78 VNB N_A_1068_21#_c_1250_n 0.00849591f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.71
cc_79 VNB N_A_1068_21#_c_1251_n 0.0475952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1068_21#_c_1252_n 0.00403568f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_81 VNB N_A_1068_21#_c_1253_n 9.88443e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1068_21#_c_1254_n 0.0160032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_887_139#_M1038_g 0.0470509f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_84 VNB N_A_887_139#_M1040_g 0.0292655f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_85 VNB N_A_887_139#_c_1345_n 0.0072322f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_86 VNB N_A_887_139#_c_1346_n 0.00950674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_887_139#_c_1347_n 0.00619557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1972_99#_M1046_g 0.0263821f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_89 VNB N_A_1972_99#_c_1474_n 0.00758877f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.71
cc_90 VNB N_A_1972_99#_c_1475_n 0.00872514f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.875
cc_91 VNB N_A_1972_99#_M1006_g 0.0282678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1972_99#_c_1477_n 0.031871f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_93 VNB N_A_1972_99#_c_1478_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1972_99#_c_1479_n 0.0203484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1972_99#_c_1480_n 0.00403324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1972_99#_c_1481_n 0.0175898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1972_99#_c_1482_n 0.00104802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1972_99#_c_1483_n 0.00911421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1972_99#_c_1484_n 0.0377313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1972_99#_c_1485_n 0.00578264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2216_99#_c_1616_n 0.017515f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.725
cc_102 VNB N_A_2216_99#_c_1617_n 0.0103367f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.71
cc_103 VNB N_A_2216_99#_c_1618_n 0.0230638f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.875
cc_104 VNB N_A_2216_99#_M1024_g 0.019445f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_105 VNB N_A_2216_99#_c_1620_n 0.0297603f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_106 VNB N_A_2216_99#_c_1621_n 0.0104651f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_107 VNB N_A_2216_99#_c_1622_n 0.0397279f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.54
cc_108 VNB N_A_2216_99#_c_1623_n 0.00360858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2216_99#_c_1624_n 0.0255844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2216_99#_c_1625_n 0.00177503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2216_99#_c_1626_n 0.0215399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2216_99#_c_1627_n 5.68909e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2216_99#_c_1628_n 0.00749017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2216_99#_c_1629_n 4.45556e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2216_99#_c_1630_n 0.0246897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2216_99#_c_1631_n 0.00690561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2216_99#_c_1632_n 0.00322117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2216_99#_c_1633_n 0.0486814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2216_99#_c_1634_n 0.0289007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1728_125#_M1051_g 0.0414372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_1728_125#_M1041_g 0.0419433f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.54
cc_122 VNB N_A_1728_125#_c_1784_n 0.0346245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_1728_125#_c_1785_n 0.0333864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1728_125#_c_1786_n 0.0119803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_1728_125#_M1007_g 0.0230856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_1728_125#_c_1788_n 0.00787249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1728_125#_c_1789_n 0.00713924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1728_125#_c_1790_n 0.0187621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_SET_B_M1003_g 0.0365192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_SET_B_M1027_g 0.00773753f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.725
cc_131 VNB N_SET_B_c_2001_n 0.252706f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_132 VNB N_SET_B_c_2002_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.205
cc_133 VNB N_SET_B_M1008_g 0.0329376f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_134 VNB N_SET_B_c_2004_n 0.247499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_SET_B_c_2005_n 0.0210256f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.54
cc_136 VNB N_SET_B_c_2006_n 0.00779893f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_137 VNB N_SET_B_c_2007_n 0.058994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_SET_B_c_2008_n 0.0126578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_SET_B_c_2009_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB SET_B 0.00165348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_SET_B_c_2011_n 0.0102347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_SET_B_c_2012_n 0.018419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_CLK_M1015_g 0.0492187f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.805
cc_144 VNB CLK 0.00310527f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_145 VNB N_CLK_c_2123_n 0.0352838f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_146 VNB N_SLEEP_B_M1014_g 0.0173227f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.805
cc_147 VNB N_SLEEP_B_M1026_g 0.00611955f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.725
cc_148 VNB N_SLEEP_B_M1049_g 0.0178973f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.71
cc_149 VNB N_SLEEP_B_M1020_g 0.0242959f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_150 VNB N_SLEEP_B_M1022_g 0.0275422f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_151 VNB N_SLEEP_B_c_2167_n 0.00620611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_SLEEP_B_c_2168_n 0.00144669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_SLEEP_B_c_2169_n 0.106066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_3466_403#_M1004_g 0.00905318f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.37
cc_155 VNB N_A_3466_403#_c_2239_n 0.00693409f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.37
cc_156 VNB N_A_3466_403#_c_2240_n 0.0109216f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.54
cc_157 VNB N_A_3466_403#_c_2241_n 0.0404865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_A_3466_403#_c_2242_n 0.00621596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_A_3466_403#_c_2243_n 0.00294342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_A_3466_403#_c_2244_n 0.00528502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_A_3466_403#_c_2245_n 0.0207142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VPWR_c_2354_n 0.780656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_A_189_119#_c_2519_n 0.00586786f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_164 VNB N_A_189_119#_c_2520_n 0.00522105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_A_189_119#_c_2521_n 0.00789731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_A_189_119#_c_2522_n 0.00291629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_A_189_119#_c_2523_n 0.00489268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_A_189_119#_c_2524_n 0.0097669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_A_189_119#_c_2525_n 0.00573585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_A_1541_125#_c_2636_n 0.0017535f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.37
cc_171 VNB N_A_1541_125#_c_2637_n 8.58533e-19 $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_172 VNB N_Q_c_2818_n 0.061358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2832_n 0.0117383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2833_n 0.043674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2834_n 0.0222572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2835_n 0.00803595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2836_n 0.0059468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2837_n 0.00517455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2838_n 0.0106025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2839_n 0.0195828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2840_n 0.0183912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2841_n 0.00494072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2842_n 0.00591524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2843_n 0.0452959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2844_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2845_n 0.0314629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2846_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2847_n 0.0933017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_VGND_c_2848_n 0.00453961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_VGND_c_2849_n 0.0196163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_191 VNB N_VGND_c_2850_n 0.051492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_192 VNB N_VGND_c_2851_n 0.08001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_193 VNB N_VGND_c_2852_n 0.0423819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_194 VNB N_VGND_c_2853_n 0.015582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_195 VNB N_VGND_c_2854_n 0.885868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_196 VNB N_VGND_c_2855_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_197 VNB N_VGND_c_2856_n 0.00510363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_198 VNB N_VGND_c_2857_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_199 VNB N_VGND_c_2858_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_200 VNB N_VGND_c_2859_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_201 VNB N_A_2074_125#_c_3022_n 0.00513591f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.37
cc_202 VNB N_A_2074_125#_c_3023_n 0.0154997f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.71
cc_203 VNB N_A_2074_125#_c_3024_n 0.00296373f $X=-0.19 $Y=-0.245 $X2=0.39
+ $Y2=1.875
cc_204 VNB N_A_2074_125#_c_3025_n 0.0052748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_205 VPB N_SCD_M1000_g 0.0492442f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.725
cc_206 VPB N_SCD_c_360_n 0.00398445f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.71
cc_207 VPB N_SCD_c_365_n 0.0168098f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.875
cc_208 VPB SCD 0.0118804f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_209 VPB N_D_M1012_g 0.0381968f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.725
cc_210 VPB N_D_c_395_n 0.0216226f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.875
cc_211 VPB N_D_c_396_n 0.00187574f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_212 VPB N_A_339_93#_M1048_g 0.0409386f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_213 VPB N_A_339_93#_c_435_n 0.0123948f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_214 VPB N_A_339_93#_c_436_n 0.0426911f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_215 VPB N_SCE_c_483_n 0.0204158f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.805
cc_216 VPB N_SCE_M1042_g 0.0194914f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_217 VPB N_SCE_M1036_g 0.0327296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_SCE_c_495_n 0.0172795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_689_139#_c_589_n 0.0616983f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_220 VPB N_A_689_139#_c_590_n 0.0182993f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.205
cc_221 VPB N_A_689_139#_M1005_g 0.0291501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_689_139#_M1021_g 0.0247893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_689_139#_c_571_n 0.00883841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_689_139#_c_574_n 0.0023433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_689_139#_c_576_n 0.0125353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_689_139#_c_596_n 0.00563237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_689_139#_c_597_n 0.0111978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_689_139#_c_598_n 0.0457462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_689_139#_c_599_n 0.00349174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_689_139#_c_600_n 0.00509541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_689_139#_c_601_n 0.00231395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_689_139#_c_602_n 0.0071901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_689_139#_c_603_n 0.0484026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_689_139#_c_580_n 0.0050676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_689_139#_c_581_n 9.56173e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_689_139#_c_582_n 6.55978e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_689_139#_c_583_n 0.0277426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_689_139#_c_585_n 0.00230456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_689_139#_c_609_n 0.00311191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_689_139#_c_610_n 9.22715e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_689_139#_c_586_n 0.00632465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_689_139#_c_587_n 0.016407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_659_113#_c_897_n 0.0556121f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.205
cc_244 VPB N_A_659_113#_M1034_g 0.0695764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_659_113#_c_930_n 0.0178299f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.54
cc_246 VPB N_A_659_113#_c_931_n 0.00719891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_659_113#_c_932_n 0.00965296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_659_113#_c_933_n 0.0186153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_659_113#_c_934_n 0.0461103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_659_113#_M1050_g 0.0232641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_659_113#_c_936_n 0.0323617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_659_113#_c_937_n 0.00922895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_659_113#_c_938_n 0.00655075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_659_113#_c_939_n 0.00476841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_659_113#_c_940_n 0.0351313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_659_113#_c_919_n 0.0209754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_659_113#_c_925_n 0.00222707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_659_113#_c_926_n 0.00153816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_659_113#_c_944_n 0.00460302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_1068_21#_M1035_g 0.0196627f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_261 VPB N_A_1068_21#_c_1256_n 0.00596691f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.54
cc_262 VPB N_A_1068_21#_c_1257_n 0.0289887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_1068_21#_c_1258_n 0.00218234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_1068_21#_c_1259_n 0.00300755f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_1068_21#_c_1254_n 0.027745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_887_139#_M1009_g 0.0443411f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_267 VPB N_A_887_139#_M1038_g 0.00609341f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_268 VPB N_A_887_139#_M1032_g 0.0250684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_887_139#_c_1345_n 0.00643902f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.54
cc_270 VPB N_A_887_139#_c_1352_n 0.00612289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_887_139#_c_1353_n 0.00374465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_887_139#_c_1354_n 0.00273658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_887_139#_c_1355_n 0.00132265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_887_139#_c_1356_n 0.0278671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_887_139#_c_1357_n 0.00858855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_887_139#_c_1346_n 0.0388113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_887_139#_c_1359_n 0.00305291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_887_139#_c_1360_n 0.0130222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_1972_99#_c_1486_n 0.0312336f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.54
cc_280 VPB N_A_1972_99#_c_1479_n 0.0174402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_A_1972_99#_c_1488_n 0.0060931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_A_1972_99#_c_1489_n 0.0100185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_1972_99#_c_1480_n 0.0052511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_1972_99#_c_1491_n 0.00455715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_A_1972_99#_c_1492_n 0.0390984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_A_1972_99#_c_1493_n 0.00210859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_A_1972_99#_c_1485_n 0.015365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_A_2216_99#_M1024_g 0.0441403f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_289 VPB N_A_2216_99#_c_1631_n 0.00553531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_A_1728_125#_c_1791_n 0.0645262f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.71
cc_291 VPB N_A_1728_125#_c_1792_n 0.0492363f $X=-0.19 $Y=1.655 $X2=0.39
+ $Y2=1.875
cc_292 VPB N_A_1728_125#_c_1793_n 0.00976808f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_293 VPB N_A_1728_125#_M1051_g 0.00554486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_A_1728_125#_c_1795_n 0.0269605f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_295 VPB N_A_1728_125#_M1041_g 0.00406f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.54
cc_296 VPB N_A_1728_125#_c_1797_n 0.0337659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_A_1728_125#_c_1798_n 0.021109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_A_1728_125#_c_1799_n 0.0170588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_A_1728_125#_c_1800_n 7.70999e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_A_1728_125#_c_1801_n 0.0486877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_A_1728_125#_c_1802_n 0.0150452f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_A_1728_125#_c_1803_n 0.00911501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_A_1728_125#_c_1788_n 0.00816475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_A_1728_125#_c_1805_n 4.40444e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_A_1728_125#_c_1789_n 5.50081e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_A_1728_125#_c_1790_n 0.0262064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_A_1728_125#_c_1808_n 0.0484092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_SET_B_M1027_g 0.0404001f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.725
cc_309 VPB N_SET_B_M1043_g 0.0240185f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_310 VPB N_SET_B_c_2011_n 0.0200526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_CLK_M1039_g 0.0264719f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.725
cc_312 VPB CLK 0.00444994f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_313 VPB N_CLK_c_2123_n 0.0119965f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.54
cc_314 VPB N_SLEEP_B_M1026_g 0.0274024f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.725
cc_315 VPB N_SLEEP_B_c_2171_n 0.036072f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_316 VPB N_SLEEP_B_c_2167_n 0.00799633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_317 VPB N_SLEEP_B_c_2168_n 0.00578675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_318 VPB N_A_3466_403#_M1004_g 0.0262963f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_319 VPB N_A_3466_403#_c_2247_n 0.00142653f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.58
cc_320 VPB N_A_3466_403#_c_2248_n 0.00268069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_321 VPB N_A_3466_403#_c_2243_n 0.00314679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_A_27_481#_c_2300_n 0.0290697f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_323 VPB N_A_27_481#_c_2301_n 0.0123991f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.71
cc_324 VPB N_A_27_481#_c_2302_n 0.0107304f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.875
cc_325 VPB N_A_27_481#_c_2303_n 0.00124656f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_326 VPB N_A_27_481#_c_2304_n 0.0111187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_A_27_481#_c_2305_n 9.09959e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_A_27_481#_c_2306_n 0.00758811f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_329 VPB N_VPWR_c_2355_n 0.00872237f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_330 VPB N_VPWR_c_2356_n 0.0315008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2357_n 0.00529899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_2358_n 0.00881296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_2359_n 0.0162187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2360_n 0.0743451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_2361_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_2362_n 0.0182105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_2363_n 0.0544409f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_338 VPB N_VPWR_c_2364_n 0.0269569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_2365_n 0.253611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_2366_n 0.0157411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_2354_n 0.104206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_342 VPB N_VPWR_c_2368_n 0.0047791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_2369_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_2370_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_2371_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_346 VPB N_A_189_119#_c_2526_n 0.0118121f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_347 VPB N_A_189_119#_c_2527_n 0.00585174f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.54
cc_348 VPB N_A_189_119#_c_2528_n 0.0141344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_349 VPB N_A_189_119#_c_2529_n 0.00349359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_350 VPB N_A_189_119#_c_2523_n 0.0381106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_351 VPB N_A_189_119#_c_2531_n 0.00570225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_352 VPB N_A_189_119#_c_2525_n 0.0043534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_353 VPB N_A_1541_125#_c_2637_n 0.00947807f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_354 VPB N_KAPWR_c_2675_n 0.00726573f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.205
cc_355 VPB N_KAPWR_c_2676_n 0.00604957f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_356 VPB N_KAPWR_c_2677_n 0.0977283f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_357 VPB N_KAPWR_c_2678_n 0.0116991f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.54
cc_358 VPB N_Q_c_2818_n 0.0501121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_359 SCD N_D_M1016_g 0.0017383f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_360 SCD N_D_c_395_n 3.38011e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_361 SCD N_D_c_396_n 0.0208019f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_362 SCD N_SCE_c_483_n 0.0176482f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_363 N_SCD_c_362_n N_SCE_c_483_n 0.02396f $X=0.39 $Y=1.37 $X2=0 $Y2=0
cc_364 N_SCD_M1001_g N_SCE_M1013_g 0.0333964f $X=0.48 $Y=0.805 $X2=0 $Y2=0
cc_365 N_SCD_M1000_g N_SCE_M1042_g 0.0189049f $X=0.48 $Y=2.725 $X2=0 $Y2=0
cc_366 N_SCD_M1001_g N_SCE_c_489_n 0.02396f $X=0.48 $Y=0.805 $X2=0 $Y2=0
cc_367 SCD N_SCE_c_489_n 0.00566255f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_368 N_SCD_c_365_n N_SCE_c_495_n 0.02396f $X=0.39 $Y=1.875 $X2=0 $Y2=0
cc_369 N_SCD_M1000_g N_A_27_481#_c_2300_n 0.0136062f $X=0.48 $Y=2.725 $X2=0
+ $Y2=0
cc_370 N_SCD_M1000_g N_A_27_481#_c_2301_n 0.00780083f $X=0.48 $Y=2.725 $X2=0
+ $Y2=0
cc_371 SCD N_A_27_481#_c_2301_n 0.0323648f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_372 N_SCD_M1000_g N_A_27_481#_c_2302_n 0.00419718f $X=0.48 $Y=2.725 $X2=0
+ $Y2=0
cc_373 N_SCD_c_365_n N_A_27_481#_c_2302_n 0.00483226f $X=0.39 $Y=1.875 $X2=0
+ $Y2=0
cc_374 SCD N_A_27_481#_c_2302_n 0.0273771f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_375 N_SCD_M1000_g N_A_27_481#_c_2303_n 7.14215e-19 $X=0.48 $Y=2.725 $X2=0
+ $Y2=0
cc_376 N_SCD_M1000_g N_VPWR_c_2355_n 0.00646225f $X=0.48 $Y=2.725 $X2=0 $Y2=0
cc_377 N_SCD_M1000_g N_VPWR_c_2362_n 0.00502664f $X=0.48 $Y=2.725 $X2=0 $Y2=0
cc_378 N_SCD_M1000_g N_VPWR_c_2354_n 0.00539301f $X=0.48 $Y=2.725 $X2=0 $Y2=0
cc_379 N_SCD_M1001_g N_A_189_119#_c_2524_n 0.00130204f $X=0.48 $Y=0.805 $X2=0
+ $Y2=0
cc_380 N_SCD_M1000_g N_KAPWR_c_2677_n 0.00451839f $X=0.48 $Y=2.725 $X2=0 $Y2=0
cc_381 N_SCD_M1001_g N_VGND_c_2833_n 0.0141223f $X=0.48 $Y=0.805 $X2=0 $Y2=0
cc_382 SCD N_VGND_c_2833_n 0.027293f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_383 N_SCD_c_362_n N_VGND_c_2833_n 0.00483226f $X=0.39 $Y=1.37 $X2=0 $Y2=0
cc_384 N_SCD_M1001_g N_VGND_c_2843_n 0.0035863f $X=0.48 $Y=0.805 $X2=0 $Y2=0
cc_385 N_SCD_M1001_g N_VGND_c_2854_n 0.00401353f $X=0.48 $Y=0.805 $X2=0 $Y2=0
cc_386 N_D_M1016_g N_A_339_93#_M1023_g 0.0387434f $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_387 N_D_M1012_g N_A_339_93#_M1048_g 0.0364183f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_388 N_D_c_395_n N_A_339_93#_c_436_n 0.0223288f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_389 N_D_c_396_n N_A_339_93#_c_436_n 3.30722e-19 $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_390 N_D_M1016_g N_SCE_c_483_n 0.0100674f $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_391 N_D_M1012_g N_SCE_c_483_n 0.00670282f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_392 N_D_c_395_n N_SCE_c_483_n 0.0195298f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_393 N_D_c_396_n N_SCE_c_483_n 0.00204407f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_394 N_D_M1016_g N_SCE_M1013_g 0.0198937f $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_395 N_D_M1016_g N_SCE_c_485_n 0.0100166f $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_396 N_D_M1012_g N_SCE_c_495_n 0.0573795f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_397 N_D_M1012_g N_A_27_481#_c_2301_n 0.00188598f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_398 N_D_c_395_n N_A_27_481#_c_2301_n 0.00151422f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_399 N_D_c_396_n N_A_27_481#_c_2301_n 0.00902013f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_400 N_D_M1012_g N_A_27_481#_c_2303_n 0.00637081f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_401 N_D_M1012_g N_A_27_481#_c_2304_n 0.010364f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_402 N_D_M1012_g N_VPWR_c_2363_n 0.00325902f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_403 N_D_M1012_g N_VPWR_c_2354_n 0.00423331f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_404 N_D_M1016_g N_A_189_119#_c_2519_n 0.0101744f $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_405 N_D_c_395_n N_A_189_119#_c_2519_n 0.00183186f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_406 N_D_c_396_n N_A_189_119#_c_2519_n 0.00544905f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_407 N_D_M1016_g N_A_189_119#_c_2524_n 0.00811291f $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_408 N_D_c_395_n N_A_189_119#_c_2524_n 0.00181663f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_409 N_D_c_396_n N_A_189_119#_c_2524_n 0.00593688f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_410 N_D_M1012_g N_A_189_119#_c_2531_n 0.00918006f $X=1.38 $Y=2.725 $X2=0
+ $Y2=0
cc_411 N_D_M1016_g N_A_189_119#_c_2525_n 0.0100412f $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_412 N_D_c_395_n N_A_189_119#_c_2525_n 0.00710199f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_413 N_D_c_396_n N_A_189_119#_c_2525_n 0.0248561f $X=1.29 $Y=1.71 $X2=0 $Y2=0
cc_414 N_D_M1012_g N_KAPWR_c_2677_n 0.00761156f $X=1.38 $Y=2.725 $X2=0 $Y2=0
cc_415 N_D_M1016_g N_VGND_c_2854_n 9.39239e-19 $X=1.3 $Y=0.805 $X2=0 $Y2=0
cc_416 N_A_339_93#_M1023_g N_SCE_c_485_n 0.0102456f $X=1.77 $Y=0.805 $X2=0 $Y2=0
cc_417 N_A_339_93#_c_437_n N_SCE_c_485_n 0.00570631f $X=2.655 $Y=0.84 $X2=0
+ $Y2=0
cc_418 N_A_339_93#_c_435_n N_SCE_M1036_g 0.0181102f $X=2.1 $Y=1.47 $X2=0 $Y2=0
cc_419 N_A_339_93#_c_434_n N_SCE_M1029_g 0.00529514f $X=2.47 $Y=1.305 $X2=0
+ $Y2=0
cc_420 N_A_339_93#_c_437_n N_SCE_M1029_g 4.26663e-19 $X=2.655 $Y=0.84 $X2=0
+ $Y2=0
cc_421 N_A_339_93#_c_434_n SCE 0.00983983f $X=2.47 $Y=1.305 $X2=0 $Y2=0
cc_422 N_A_339_93#_c_435_n SCE 0.0215723f $X=2.1 $Y=1.47 $X2=0 $Y2=0
cc_423 N_A_339_93#_c_437_n SCE 0.00115924f $X=2.655 $Y=0.84 $X2=0 $Y2=0
cc_424 N_A_339_93#_c_434_n N_SCE_c_491_n 0.00188817f $X=2.47 $Y=1.305 $X2=0
+ $Y2=0
cc_425 N_A_339_93#_c_435_n N_SCE_c_491_n 0.00733591f $X=2.1 $Y=1.47 $X2=0 $Y2=0
cc_426 N_A_339_93#_c_436_n N_SCE_c_491_n 0.0135432f $X=2.1 $Y=1.47 $X2=0 $Y2=0
cc_427 N_A_339_93#_c_437_n N_SCE_c_491_n 0.00136269f $X=2.655 $Y=0.84 $X2=0
+ $Y2=0
cc_428 N_A_339_93#_M1048_g N_A_27_481#_c_2304_n 0.00901726f $X=1.81 $Y=2.725
+ $X2=0 $Y2=0
cc_429 N_A_339_93#_M1048_g N_A_27_481#_c_2306_n 0.00260904f $X=1.81 $Y=2.725
+ $X2=0 $Y2=0
cc_430 N_A_339_93#_M1048_g N_VPWR_c_2363_n 0.00325902f $X=1.81 $Y=2.725 $X2=0
+ $Y2=0
cc_431 N_A_339_93#_M1048_g N_VPWR_c_2354_n 0.00518531f $X=1.81 $Y=2.725 $X2=0
+ $Y2=0
cc_432 N_A_339_93#_M1023_g N_A_189_119#_c_2519_n 0.00552172f $X=1.77 $Y=0.805
+ $X2=0 $Y2=0
cc_433 N_A_339_93#_M1036_s N_A_189_119#_c_2526_n 0.00620515f $X=2.425 $Y=1.795
+ $X2=0 $Y2=0
cc_434 N_A_339_93#_M1048_g N_A_189_119#_c_2526_n 0.0141445f $X=1.81 $Y=2.725
+ $X2=0 $Y2=0
cc_435 N_A_339_93#_c_435_n N_A_189_119#_c_2526_n 0.0582121f $X=2.1 $Y=1.47 $X2=0
+ $Y2=0
cc_436 N_A_339_93#_c_436_n N_A_189_119#_c_2526_n 0.00390699f $X=2.1 $Y=1.47
+ $X2=0 $Y2=0
cc_437 N_A_339_93#_M1023_g N_A_189_119#_c_2524_n 0.0014734f $X=1.77 $Y=0.805
+ $X2=0 $Y2=0
cc_438 N_A_339_93#_M1048_g N_A_189_119#_c_2531_n 0.0126776f $X=1.81 $Y=2.725
+ $X2=0 $Y2=0
cc_439 N_A_339_93#_M1023_g N_A_189_119#_c_2525_n 0.00847653f $X=1.77 $Y=0.805
+ $X2=0 $Y2=0
cc_440 N_A_339_93#_M1048_g N_A_189_119#_c_2525_n 0.00960126f $X=1.81 $Y=2.725
+ $X2=0 $Y2=0
cc_441 N_A_339_93#_c_434_n N_A_189_119#_c_2525_n 0.00726118f $X=2.47 $Y=1.305
+ $X2=0 $Y2=0
cc_442 N_A_339_93#_c_435_n N_A_189_119#_c_2525_n 0.0571887f $X=2.1 $Y=1.47 $X2=0
+ $Y2=0
cc_443 N_A_339_93#_c_436_n N_A_189_119#_c_2525_n 0.0185823f $X=2.1 $Y=1.47 $X2=0
+ $Y2=0
cc_444 N_A_339_93#_M1048_g N_KAPWR_c_2677_n 0.00192067f $X=1.81 $Y=2.725 $X2=0
+ $Y2=0
cc_445 N_A_339_93#_M1023_g N_VGND_c_2834_n 0.0119963f $X=1.77 $Y=0.805 $X2=0
+ $Y2=0
cc_446 N_A_339_93#_c_434_n N_VGND_c_2834_n 0.00176105f $X=2.47 $Y=1.305 $X2=0
+ $Y2=0
cc_447 N_A_339_93#_c_435_n N_VGND_c_2834_n 0.0156175f $X=2.1 $Y=1.47 $X2=0 $Y2=0
cc_448 N_A_339_93#_c_436_n N_VGND_c_2834_n 0.00183955f $X=2.1 $Y=1.47 $X2=0
+ $Y2=0
cc_449 N_A_339_93#_c_437_n N_VGND_c_2834_n 0.024902f $X=2.655 $Y=0.84 $X2=0
+ $Y2=0
cc_450 N_A_339_93#_c_437_n N_VGND_c_2835_n 0.0127193f $X=2.655 $Y=0.84 $X2=0
+ $Y2=0
cc_451 N_A_339_93#_c_437_n N_VGND_c_2849_n 0.00625484f $X=2.655 $Y=0.84 $X2=0
+ $Y2=0
cc_452 N_A_339_93#_M1023_g N_VGND_c_2854_n 9.39239e-19 $X=1.77 $Y=0.805 $X2=0
+ $Y2=0
cc_453 N_A_339_93#_c_437_n N_VGND_c_2854_n 0.00872741f $X=2.655 $Y=0.84 $X2=0
+ $Y2=0
cc_454 N_SCE_M1036_g N_A_689_139#_c_571_n 0.0027751f $X=2.77 $Y=2.115 $X2=0
+ $Y2=0
cc_455 N_SCE_M1029_g N_A_689_139#_c_571_n 9.3167e-19 $X=2.87 $Y=0.905 $X2=0
+ $Y2=0
cc_456 SCE N_A_689_139#_c_571_n 0.0295304f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_457 N_SCE_c_491_n N_A_689_139#_c_571_n 5.69415e-19 $X=2.89 $Y=1.39 $X2=0
+ $Y2=0
cc_458 N_SCE_M1029_g N_A_689_139#_c_579_n 0.00128934f $X=2.87 $Y=0.905 $X2=0
+ $Y2=0
cc_459 N_SCE_M1036_g N_A_689_139#_c_602_n 0.00209451f $X=2.77 $Y=2.115 $X2=0
+ $Y2=0
cc_460 N_SCE_M1029_g N_A_659_113#_c_896_n 0.0148512f $X=2.87 $Y=0.905 $X2=0
+ $Y2=0
cc_461 SCE N_A_659_113#_c_896_n 0.00173869f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_462 N_SCE_M1036_g N_A_659_113#_c_897_n 0.0189367f $X=2.77 $Y=2.115 $X2=0
+ $Y2=0
cc_463 SCE N_A_659_113#_c_897_n 7.30348e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_464 N_SCE_c_491_n N_A_659_113#_c_897_n 0.00559859f $X=2.89 $Y=1.39 $X2=0
+ $Y2=0
cc_465 N_SCE_c_491_n N_A_659_113#_c_899_n 0.0082579f $X=2.89 $Y=1.39 $X2=0 $Y2=0
cc_466 N_SCE_M1042_g N_A_27_481#_c_2300_n 6.9536e-19 $X=0.99 $Y=2.725 $X2=0
+ $Y2=0
cc_467 N_SCE_c_483_n N_A_27_481#_c_2301_n 0.00584112f $X=0.84 $Y=2.085 $X2=0
+ $Y2=0
cc_468 N_SCE_c_495_n N_A_27_481#_c_2301_n 0.0115865f $X=0.99 $Y=2.16 $X2=0 $Y2=0
cc_469 N_SCE_M1042_g N_A_27_481#_c_2303_n 0.0121514f $X=0.99 $Y=2.725 $X2=0
+ $Y2=0
cc_470 N_SCE_c_495_n N_A_27_481#_c_2303_n 5.48408e-19 $X=0.99 $Y=2.16 $X2=0
+ $Y2=0
cc_471 N_SCE_M1042_g N_A_27_481#_c_2305_n 0.00390882f $X=0.99 $Y=2.725 $X2=0
+ $Y2=0
cc_472 N_SCE_M1042_g N_VPWR_c_2355_n 0.00436122f $X=0.99 $Y=2.725 $X2=0 $Y2=0
cc_473 N_SCE_c_495_n N_VPWR_c_2355_n 0.00234309f $X=0.99 $Y=2.16 $X2=0 $Y2=0
cc_474 N_SCE_M1042_g N_VPWR_c_2363_n 0.0047293f $X=0.99 $Y=2.725 $X2=0 $Y2=0
cc_475 N_SCE_M1036_g N_VPWR_c_2363_n 0.00297774f $X=2.77 $Y=2.115 $X2=0 $Y2=0
cc_476 N_SCE_M1042_g N_VPWR_c_2354_n 0.00466629f $X=0.99 $Y=2.725 $X2=0 $Y2=0
cc_477 N_SCE_c_485_n N_A_189_119#_c_2519_n 0.00645921f $X=2.795 $Y=0.18 $X2=0
+ $Y2=0
cc_478 N_SCE_M1036_g N_A_189_119#_c_2526_n 0.0159377f $X=2.77 $Y=2.115 $X2=0
+ $Y2=0
cc_479 SCE N_A_189_119#_c_2526_n 0.0125397f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_480 N_SCE_c_491_n N_A_189_119#_c_2526_n 0.00324635f $X=2.89 $Y=1.39 $X2=0
+ $Y2=0
cc_481 N_SCE_M1013_g N_A_189_119#_c_2524_n 0.0100033f $X=0.87 $Y=0.805 $X2=0
+ $Y2=0
cc_482 N_SCE_c_485_n N_A_189_119#_c_2524_n 0.00381922f $X=2.795 $Y=0.18 $X2=0
+ $Y2=0
cc_483 N_SCE_c_495_n N_A_189_119#_c_2531_n 4.79185e-19 $X=0.99 $Y=2.16 $X2=0
+ $Y2=0
cc_484 N_SCE_M1042_g N_KAPWR_c_2677_n 0.00202335f $X=0.99 $Y=2.725 $X2=0 $Y2=0
cc_485 N_SCE_M1036_g N_KAPWR_c_2677_n 0.00469573f $X=2.77 $Y=2.115 $X2=0 $Y2=0
cc_486 N_SCE_c_495_n N_KAPWR_c_2677_n 0.00169078f $X=0.99 $Y=2.16 $X2=0 $Y2=0
cc_487 N_SCE_M1013_g N_VGND_c_2833_n 0.0018473f $X=0.87 $Y=0.805 $X2=0 $Y2=0
cc_488 N_SCE_c_486_n N_VGND_c_2833_n 0.00977077f $X=0.945 $Y=0.18 $X2=0 $Y2=0
cc_489 N_SCE_c_485_n N_VGND_c_2834_n 0.0216291f $X=2.795 $Y=0.18 $X2=0 $Y2=0
cc_490 N_SCE_M1029_g N_VGND_c_2834_n 0.0100548f $X=2.87 $Y=0.905 $X2=0 $Y2=0
cc_491 N_SCE_c_485_n N_VGND_c_2835_n 0.00763335f $X=2.795 $Y=0.18 $X2=0 $Y2=0
cc_492 N_SCE_M1029_g N_VGND_c_2835_n 0.0299792f $X=2.87 $Y=0.905 $X2=0 $Y2=0
cc_493 SCE N_VGND_c_2835_n 0.0247102f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_494 N_SCE_c_491_n N_VGND_c_2835_n 6.13938e-19 $X=2.89 $Y=1.39 $X2=0 $Y2=0
cc_495 N_SCE_c_486_n N_VGND_c_2843_n 0.0375648f $X=0.945 $Y=0.18 $X2=0 $Y2=0
cc_496 N_SCE_c_485_n N_VGND_c_2849_n 0.0228563f $X=2.795 $Y=0.18 $X2=0 $Y2=0
cc_497 N_SCE_c_485_n N_VGND_c_2854_n 0.0678934f $X=2.795 $Y=0.18 $X2=0 $Y2=0
cc_498 N_SCE_c_486_n N_VGND_c_2854_n 0.0107881f $X=0.945 $Y=0.18 $X2=0 $Y2=0
cc_499 N_A_689_139#_c_571_n N_A_659_113#_c_896_n 0.0132222f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_500 N_A_689_139#_c_579_n N_A_659_113#_c_896_n 9.7247e-19 $X=4.015 $Y=0.42
+ $X2=0 $Y2=0
cc_501 N_A_689_139#_c_588_n N_A_659_113#_c_896_n 0.00110296f $X=3.85 $Y=0.18
+ $X2=0 $Y2=0
cc_502 N_A_689_139#_c_571_n N_A_659_113#_c_897_n 0.0139138f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_503 N_A_689_139#_c_601_n N_A_659_113#_c_897_n 8.68414e-19 $X=4.132 $Y=1.89
+ $X2=0 $Y2=0
cc_504 N_A_689_139#_c_602_n N_A_659_113#_c_897_n 0.0110007f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_505 N_A_689_139#_c_603_n N_A_659_113#_c_897_n 0.013438f $X=4.17 $Y=1.89 $X2=0
+ $Y2=0
cc_506 N_A_689_139#_c_571_n N_A_659_113#_c_898_n 0.0123675f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_507 N_A_689_139#_c_579_n N_A_659_113#_c_898_n 0.00118168f $X=4.015 $Y=0.42
+ $X2=0 $Y2=0
cc_508 N_A_689_139#_c_602_n N_A_659_113#_c_898_n 0.007979f $X=4.17 $Y=1.89 $X2=0
+ $Y2=0
cc_509 N_A_689_139#_c_603_n N_A_659_113#_c_898_n 0.0108462f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_510 N_A_689_139#_c_588_n N_A_659_113#_c_898_n 0.0060778f $X=3.85 $Y=0.18
+ $X2=0 $Y2=0
cc_511 N_A_689_139#_c_571_n N_A_659_113#_c_899_n 0.00434296f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_512 N_A_689_139#_c_579_n N_A_659_113#_c_899_n 2.73184e-19 $X=4.015 $Y=0.42
+ $X2=0 $Y2=0
cc_513 N_A_689_139#_c_567_n N_A_659_113#_c_900_n 0.00518713f $X=4.83 $Y=0.18
+ $X2=0 $Y2=0
cc_514 N_A_689_139#_c_568_n N_A_659_113#_c_900_n 0.00752782f $X=4.905 $Y=0.255
+ $X2=0 $Y2=0
cc_515 N_A_689_139#_c_571_n N_A_659_113#_c_900_n 0.00432191f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_516 N_A_689_139#_c_572_n N_A_659_113#_c_900_n 0.00315349f $X=5.11 $Y=0.34
+ $X2=0 $Y2=0
cc_517 N_A_689_139#_c_573_n N_A_659_113#_c_900_n 3.65704e-19 $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_518 N_A_689_139#_c_588_n N_A_659_113#_c_900_n 8.84721e-19 $X=3.85 $Y=0.18
+ $X2=0 $Y2=0
cc_519 N_A_689_139#_c_568_n N_A_659_113#_c_901_n 0.0064846f $X=4.905 $Y=0.255
+ $X2=0 $Y2=0
cc_520 N_A_689_139#_c_573_n N_A_659_113#_c_901_n 0.0140068f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_521 N_A_689_139#_c_580_n N_A_659_113#_c_901_n 0.005786f $X=5.95 $Y=1.592
+ $X2=0 $Y2=0
cc_522 N_A_689_139#_c_589_n N_A_659_113#_M1034_g 0.0276183f $X=5.08 $Y=2.32
+ $X2=0 $Y2=0
cc_523 N_A_689_139#_c_573_n N_A_659_113#_M1034_g 0.00213586f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_524 N_A_689_139#_c_580_n N_A_659_113#_M1034_g 0.0128003f $X=5.95 $Y=1.592
+ $X2=0 $Y2=0
cc_525 N_A_689_139#_c_581_n N_A_659_113#_M1034_g 8.75187e-19 $X=6.12 $Y=1.592
+ $X2=0 $Y2=0
cc_526 N_A_689_139#_c_576_n N_A_659_113#_c_930_n 0.00298041f $X=7.93 $Y=2.905
+ $X2=0 $Y2=0
cc_527 N_A_689_139#_c_647_p N_A_659_113#_c_930_n 0.0107116f $X=8.525 $Y=2.99
+ $X2=0 $Y2=0
cc_528 N_A_689_139#_c_596_n N_A_659_113#_c_930_n 0.0140403f $X=8.61 $Y=2.905
+ $X2=0 $Y2=0
cc_529 N_A_689_139#_c_596_n N_A_659_113#_c_931_n 0.00646906f $X=8.61 $Y=2.905
+ $X2=0 $Y2=0
cc_530 N_A_689_139#_c_582_n N_A_659_113#_c_931_n 4.4451e-19 $X=8.645 $Y=1.575
+ $X2=0 $Y2=0
cc_531 N_A_689_139#_c_596_n N_A_659_113#_c_932_n 0.00208927f $X=8.61 $Y=2.905
+ $X2=0 $Y2=0
cc_532 N_A_689_139#_c_583_n N_A_659_113#_c_932_n 0.0235539f $X=8.645 $Y=1.575
+ $X2=0 $Y2=0
cc_533 N_A_689_139#_c_647_p N_A_659_113#_c_933_n 0.00132869f $X=8.525 $Y=2.99
+ $X2=0 $Y2=0
cc_534 N_A_689_139#_c_596_n N_A_659_113#_c_933_n 0.00460597f $X=8.61 $Y=2.905
+ $X2=0 $Y2=0
cc_535 N_A_689_139#_c_597_n N_A_659_113#_c_933_n 2.98852e-19 $X=9.4 $Y=2.405
+ $X2=0 $Y2=0
cc_536 N_A_689_139#_c_597_n N_A_659_113#_c_934_n 0.00434958f $X=9.4 $Y=2.405
+ $X2=0 $Y2=0
cc_537 N_A_689_139#_c_598_n N_A_659_113#_c_934_n 0.0217224f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_538 N_A_689_139#_c_609_n N_A_659_113#_c_934_n 0.00877489f $X=9.425 $Y=2.135
+ $X2=0 $Y2=0
cc_539 N_A_689_139#_c_577_n N_A_659_113#_M1050_g 0.00743921f $X=9.365 $Y=0.68
+ $X2=0 $Y2=0
cc_540 N_A_689_139#_c_583_n N_A_659_113#_M1050_g 0.0033994f $X=8.645 $Y=1.575
+ $X2=0 $Y2=0
cc_541 N_A_689_139#_c_585_n N_A_659_113#_M1050_g 0.0391081f $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_542 N_A_689_139#_c_609_n N_A_659_113#_M1050_g 0.0042145f $X=9.425 $Y=2.135
+ $X2=0 $Y2=0
cc_543 N_A_689_139#_c_609_n N_A_659_113#_c_938_n 0.00467325f $X=9.425 $Y=2.135
+ $X2=0 $Y2=0
cc_544 N_A_689_139#_c_573_n N_A_659_113#_c_905_n 0.0401002f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_545 N_A_689_139#_c_580_n N_A_659_113#_c_905_n 0.025711f $X=5.95 $Y=1.592
+ $X2=0 $Y2=0
cc_546 N_A_689_139#_c_573_n N_A_659_113#_c_906_n 0.00524736f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_547 N_A_689_139#_c_580_n N_A_659_113#_c_906_n 0.00446668f $X=5.95 $Y=1.592
+ $X2=0 $Y2=0
cc_548 N_A_689_139#_c_581_n N_A_659_113#_c_907_n 0.00113811f $X=6.12 $Y=1.592
+ $X2=0 $Y2=0
cc_549 N_A_689_139#_c_573_n N_A_659_113#_c_908_n 0.0135498f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_550 N_A_689_139#_c_575_n N_A_659_113#_c_913_n 0.0598001f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_551 N_A_689_139#_c_575_n N_A_659_113#_c_914_n 0.0143582f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_552 N_A_689_139#_M1025_g N_A_659_113#_c_915_n 7.2386e-19 $X=8.205 $Y=0.945
+ $X2=0 $Y2=0
cc_553 N_A_689_139#_M1025_g N_A_659_113#_c_916_n 0.00196625f $X=8.205 $Y=0.945
+ $X2=0 $Y2=0
cc_554 N_A_689_139#_M1017_g N_A_659_113#_c_916_n 0.00174767f $X=8.565 $Y=0.945
+ $X2=0 $Y2=0
cc_555 N_A_689_139#_c_577_n N_A_659_113#_c_916_n 0.060697f $X=9.365 $Y=0.68
+ $X2=0 $Y2=0
cc_556 N_A_689_139#_c_578_n N_A_659_113#_c_916_n 0.0129683f $X=8.695 $Y=0.68
+ $X2=0 $Y2=0
cc_557 N_A_689_139#_c_577_n N_A_659_113#_c_918_n 0.00532719f $X=9.365 $Y=0.68
+ $X2=0 $Y2=0
cc_558 N_A_689_139#_c_585_n N_A_659_113#_c_918_n 0.0220729f $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_559 N_A_689_139#_c_598_n N_A_659_113#_c_939_n 0.0131038f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_560 N_A_689_139#_c_585_n N_A_659_113#_c_939_n 0.0103436f $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_561 N_A_689_139#_c_598_n N_A_659_113#_c_940_n 0.00159887f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_562 N_A_689_139#_c_585_n N_A_659_113#_c_940_n 6.55449e-19 $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_563 N_A_689_139#_c_585_n N_A_659_113#_c_926_n 0.0055599f $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_564 N_A_689_139#_c_567_n N_A_1068_21#_c_1248_n 0.0115184f $X=4.83 $Y=0.18
+ $X2=0 $Y2=0
cc_565 N_A_689_139#_c_572_n N_A_1068_21#_c_1248_n 0.00158383f $X=5.11 $Y=0.34
+ $X2=0 $Y2=0
cc_566 N_A_689_139#_c_573_n N_A_1068_21#_c_1248_n 0.00708175f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_567 N_A_689_139#_c_580_n N_A_1068_21#_c_1249_n 0.00366135f $X=5.95 $Y=1.592
+ $X2=0 $Y2=0
cc_568 N_A_689_139#_c_581_n N_A_1068_21#_c_1249_n 5.93034e-19 $X=6.12 $Y=1.592
+ $X2=0 $Y2=0
cc_569 N_A_689_139#_c_568_n N_A_1068_21#_c_1250_n 0.0115184f $X=4.905 $Y=0.255
+ $X2=0 $Y2=0
cc_570 N_A_689_139#_c_575_n N_A_1068_21#_c_1251_n 0.00212746f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_571 N_A_689_139#_c_581_n N_A_1068_21#_c_1251_n 0.00240906f $X=6.12 $Y=1.592
+ $X2=0 $Y2=0
cc_572 N_A_689_139#_c_575_n N_A_1068_21#_c_1252_n 0.0209018f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_573 N_A_689_139#_c_581_n N_A_1068_21#_c_1252_n 0.0230505f $X=6.12 $Y=1.592
+ $X2=0 $Y2=0
cc_574 N_A_689_139#_c_575_n N_A_1068_21#_c_1254_n 0.00718514f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_575 N_A_689_139#_c_581_n N_A_1068_21#_c_1254_n 0.00674944f $X=6.12 $Y=1.592
+ $X2=0 $Y2=0
cc_576 N_A_689_139#_c_572_n N_A_887_139#_M1047_d 0.0028305f $X=5.11 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_577 N_A_689_139#_c_575_n N_A_887_139#_M1038_g 0.0144342f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_578 N_A_689_139#_c_581_n N_A_887_139#_M1038_g 3.64568e-19 $X=6.12 $Y=1.592
+ $X2=0 $Y2=0
cc_579 N_A_689_139#_M1025_g N_A_887_139#_M1040_g 0.0113367f $X=8.205 $Y=0.945
+ $X2=0 $Y2=0
cc_580 N_A_689_139#_c_575_n N_A_887_139#_M1040_g 0.00780932f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_581 N_A_689_139#_c_701_p N_A_887_139#_M1032_g 0.00153968f $X=8.015 $Y=2.99
+ $X2=0 $Y2=0
cc_582 N_A_689_139#_c_573_n N_A_887_139#_c_1345_n 0.0297075f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_583 N_A_689_139#_c_574_n N_A_887_139#_c_1345_n 0.0143582f $X=5.28 $Y=1.63
+ $X2=0 $Y2=0
cc_584 N_A_689_139#_c_589_n N_A_887_139#_c_1352_n 0.00889774f $X=5.08 $Y=2.32
+ $X2=0 $Y2=0
cc_585 N_A_689_139#_c_574_n N_A_887_139#_c_1352_n 0.00738142f $X=5.28 $Y=1.63
+ $X2=0 $Y2=0
cc_586 N_A_689_139#_c_589_n N_A_887_139#_c_1353_n 0.00436548f $X=5.08 $Y=2.32
+ $X2=0 $Y2=0
cc_587 N_A_689_139#_c_589_n N_A_887_139#_c_1354_n 0.00685819f $X=5.08 $Y=2.32
+ $X2=0 $Y2=0
cc_588 N_A_689_139#_M1005_g N_A_887_139#_c_1354_n 0.0125538f $X=5.155 $Y=2.885
+ $X2=0 $Y2=0
cc_589 N_A_689_139#_c_575_n N_A_887_139#_c_1355_n 0.0911134f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_590 N_A_689_139#_c_575_n N_A_887_139#_c_1356_n 0.00462763f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_591 N_A_689_139#_c_576_n N_A_887_139#_c_1357_n 0.0226153f $X=7.93 $Y=2.905
+ $X2=0 $Y2=0
cc_592 N_A_689_139#_c_575_n N_A_887_139#_c_1346_n 0.0113375f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_593 N_A_689_139#_c_576_n N_A_887_139#_c_1346_n 0.0216346f $X=7.93 $Y=2.905
+ $X2=0 $Y2=0
cc_594 N_A_689_139#_c_583_n N_A_887_139#_c_1346_n 0.0113367f $X=8.645 $Y=1.575
+ $X2=0 $Y2=0
cc_595 N_A_689_139#_c_568_n N_A_887_139#_c_1347_n 0.0104038f $X=4.905 $Y=0.255
+ $X2=0 $Y2=0
cc_596 N_A_689_139#_c_571_n N_A_887_139#_c_1347_n 0.00230419f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_597 N_A_689_139#_c_572_n N_A_887_139#_c_1347_n 0.0248746f $X=5.11 $Y=0.34
+ $X2=0 $Y2=0
cc_598 N_A_689_139#_c_573_n N_A_887_139#_c_1347_n 0.0367022f $X=5.195 $Y=1.545
+ $X2=0 $Y2=0
cc_599 N_A_689_139#_c_574_n N_A_887_139#_c_1359_n 0.00649231f $X=5.28 $Y=1.63
+ $X2=0 $Y2=0
cc_600 N_A_689_139#_c_580_n N_A_887_139#_c_1359_n 0.0196617f $X=5.95 $Y=1.592
+ $X2=0 $Y2=0
cc_601 N_A_689_139#_c_575_n N_A_887_139#_c_1360_n 0.0167908f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_602 N_A_689_139#_c_580_n N_A_887_139#_c_1360_n 0.0397407f $X=5.95 $Y=1.592
+ $X2=0 $Y2=0
cc_603 N_A_689_139#_c_598_n N_A_1972_99#_M1018_s 0.0140243f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_604 N_A_689_139#_c_724_p N_A_1972_99#_M1018_s 0.00412049f $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_605 N_A_689_139#_c_725_p N_A_1972_99#_M1018_s 0.0123566f $X=12.06 $Y=2.31
+ $X2=0 $Y2=0
cc_606 N_A_689_139#_c_577_n N_A_1972_99#_M1046_g 4.94074e-19 $X=9.365 $Y=0.68
+ $X2=0 $Y2=0
cc_607 N_A_689_139#_c_585_n N_A_1972_99#_M1046_g 0.00250033f $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_608 N_A_689_139#_M1021_g N_A_1972_99#_c_1479_n 0.0651518f $X=14.185 $Y=2.57
+ $X2=0 $Y2=0
cc_609 N_A_689_139#_c_586_n N_A_1972_99#_c_1479_n 0.00277569f $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_610 N_A_689_139#_c_587_n N_A_1972_99#_c_1479_n 0.0198387f $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_611 N_A_689_139#_c_598_n N_A_1972_99#_c_1488_n 0.0212356f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_612 N_A_689_139#_c_598_n N_A_1972_99#_c_1489_n 0.00726212f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_613 N_A_689_139#_c_724_p N_A_1972_99#_c_1489_n 0.0538718f $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_614 N_A_689_139#_c_725_p N_A_1972_99#_c_1489_n 0.0129609f $X=12.06 $Y=2.31
+ $X2=0 $Y2=0
cc_615 N_A_689_139#_c_610_n N_A_1972_99#_c_1489_n 0.00363015f $X=13.27 $Y=2.095
+ $X2=0 $Y2=0
cc_616 N_A_689_139#_c_600_n N_A_1972_99#_c_1481_n 0.0111637f $X=14.04 $Y=2.095
+ $X2=0 $Y2=0
cc_617 N_A_689_139#_c_610_n N_A_1972_99#_c_1481_n 0.00479559f $X=13.27 $Y=2.095
+ $X2=0 $Y2=0
cc_618 N_A_689_139#_c_586_n N_A_1972_99#_c_1481_n 0.0255349f $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_619 N_A_689_139#_c_587_n N_A_1972_99#_c_1481_n 0.00160958f $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_620 N_A_689_139#_c_598_n N_A_1972_99#_c_1491_n 0.0215838f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_621 N_A_689_139#_c_598_n N_A_1972_99#_c_1492_n 0.00224424f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_622 N_A_689_139#_c_598_n N_A_1972_99#_c_1493_n 0.0242013f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_623 N_A_689_139#_c_725_p N_A_1972_99#_c_1493_n 7.64219e-19 $X=12.06 $Y=2.31
+ $X2=0 $Y2=0
cc_624 N_A_689_139#_c_600_n N_A_2216_99#_c_1618_n 5.43971e-19 $X=14.04 $Y=2.095
+ $X2=0 $Y2=0
cc_625 N_A_689_139#_c_610_n N_A_2216_99#_c_1618_n 3.44468e-19 $X=13.27 $Y=2.095
+ $X2=0 $Y2=0
cc_626 N_A_689_139#_c_724_p N_A_2216_99#_M1024_g 0.0139059f $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_627 N_A_689_139#_c_600_n N_A_2216_99#_M1024_g 2.65691e-19 $X=14.04 $Y=2.095
+ $X2=0 $Y2=0
cc_628 N_A_689_139#_c_610_n N_A_2216_99#_M1024_g 0.0136033f $X=13.27 $Y=2.095
+ $X2=0 $Y2=0
cc_629 N_A_689_139#_c_577_n N_A_1728_125#_M1017_d 0.0178533f $X=9.365 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_630 N_A_689_139#_c_585_n N_A_1728_125#_M1017_d 0.00699335f $X=9.425 $Y=1.885
+ $X2=-0.19 $Y2=-0.245
cc_631 N_A_689_139#_c_600_n N_A_1728_125#_M1043_d 0.00172391f $X=14.04 $Y=2.095
+ $X2=0 $Y2=0
cc_632 N_A_689_139#_c_598_n N_A_1728_125#_c_1791_n 0.0153298f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_633 N_A_689_139#_c_725_p N_A_1728_125#_c_1791_n 0.00408807f $X=12.06 $Y=2.31
+ $X2=0 $Y2=0
cc_634 N_A_689_139#_c_598_n N_A_1728_125#_c_1792_n 0.00195299f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_635 N_A_689_139#_c_724_p N_A_1728_125#_c_1792_n 5.42449e-19 $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_636 N_A_689_139#_c_725_p N_A_1728_125#_c_1792_n 8.6391e-19 $X=12.06 $Y=2.31
+ $X2=0 $Y2=0
cc_637 N_A_689_139#_c_724_p N_A_1728_125#_c_1795_n 0.0165643f $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_638 N_A_689_139#_c_725_p N_A_1728_125#_c_1795_n 0.00678436f $X=12.06 $Y=2.31
+ $X2=0 $Y2=0
cc_639 N_A_689_139#_c_610_n N_A_1728_125#_c_1795_n 9.06874e-19 $X=13.27 $Y=2.095
+ $X2=0 $Y2=0
cc_640 N_A_689_139#_c_724_p N_A_1728_125#_c_1799_n 2.62245e-19 $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_641 N_A_689_139#_c_596_n N_A_1728_125#_c_1800_n 0.0245136f $X=8.61 $Y=2.905
+ $X2=0 $Y2=0
cc_642 N_A_689_139#_c_597_n N_A_1728_125#_c_1800_n 0.012894f $X=9.4 $Y=2.405
+ $X2=0 $Y2=0
cc_643 N_A_689_139#_c_647_p N_A_1728_125#_c_1823_n 0.00595868f $X=8.525 $Y=2.99
+ $X2=0 $Y2=0
cc_644 N_A_689_139#_c_596_n N_A_1728_125#_c_1823_n 0.0133251f $X=8.61 $Y=2.905
+ $X2=0 $Y2=0
cc_645 N_A_689_139#_c_599_n N_A_1728_125#_c_1825_n 0.0145003f $X=9.485 $Y=2.49
+ $X2=0 $Y2=0
cc_646 N_A_689_139#_c_598_n N_A_1728_125#_c_1801_n 0.16074f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_647 N_A_689_139#_c_599_n N_A_1728_125#_c_1801_n 0.0124259f $X=9.485 $Y=2.49
+ $X2=0 $Y2=0
cc_648 N_A_689_139#_c_724_p N_A_1728_125#_c_1801_n 0.00450579f $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_649 N_A_689_139#_c_725_p N_A_1728_125#_c_1801_n 0.0112892f $X=12.06 $Y=2.31
+ $X2=0 $Y2=0
cc_650 N_A_689_139#_c_724_p N_A_1728_125#_c_1830_n 0.0383016f $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_651 N_A_689_139#_c_600_n N_A_1728_125#_c_1830_n 0.0113652f $X=14.04 $Y=2.095
+ $X2=0 $Y2=0
cc_652 N_A_689_139#_c_610_n N_A_1728_125#_c_1830_n 0.00748276f $X=13.27 $Y=2.095
+ $X2=0 $Y2=0
cc_653 N_A_689_139#_M1017_g N_A_1728_125#_c_1833_n 0.00186886f $X=8.565 $Y=0.945
+ $X2=0 $Y2=0
cc_654 N_A_689_139#_c_577_n N_A_1728_125#_c_1833_n 0.0249664f $X=9.365 $Y=0.68
+ $X2=0 $Y2=0
cc_655 N_A_689_139#_c_585_n N_A_1728_125#_c_1833_n 0.0221168f $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_656 N_A_689_139#_M1017_g N_A_1728_125#_c_1788_n 0.00108885f $X=8.565 $Y=0.945
+ $X2=0 $Y2=0
cc_657 N_A_689_139#_c_596_n N_A_1728_125#_c_1788_n 0.0289504f $X=8.61 $Y=2.905
+ $X2=0 $Y2=0
cc_658 N_A_689_139#_c_582_n N_A_1728_125#_c_1788_n 0.0241333f $X=8.645 $Y=1.575
+ $X2=0 $Y2=0
cc_659 N_A_689_139#_c_583_n N_A_1728_125#_c_1788_n 0.00445603f $X=8.645 $Y=1.575
+ $X2=0 $Y2=0
cc_660 N_A_689_139#_c_584_n N_A_1728_125#_c_1788_n 0.00993968f $X=8.64 $Y=1.41
+ $X2=0 $Y2=0
cc_661 N_A_689_139#_c_585_n N_A_1728_125#_c_1788_n 0.0358836f $X=9.425 $Y=1.885
+ $X2=0 $Y2=0
cc_662 N_A_689_139#_c_609_n N_A_1728_125#_c_1788_n 0.0210825f $X=9.425 $Y=2.135
+ $X2=0 $Y2=0
cc_663 N_A_689_139#_c_724_p N_A_1728_125#_c_1805_n 0.00931033f $X=13.185 $Y=2.31
+ $X2=0 $Y2=0
cc_664 N_A_689_139#_M1021_g N_A_1728_125#_c_1844_n 0.00831194f $X=14.185 $Y=2.57
+ $X2=0 $Y2=0
cc_665 N_A_689_139#_c_600_n N_A_1728_125#_c_1844_n 0.012473f $X=14.04 $Y=2.095
+ $X2=0 $Y2=0
cc_666 N_A_689_139#_c_586_n N_A_1728_125#_c_1844_n 0.00530387f $X=14.205
+ $Y=1.745 $X2=0 $Y2=0
cc_667 N_A_689_139#_M1021_g N_A_1728_125#_c_1847_n 0.0122275f $X=14.185 $Y=2.57
+ $X2=0 $Y2=0
cc_668 N_A_689_139#_c_586_n N_A_1728_125#_c_1847_n 0.0102108f $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_669 N_A_689_139#_M1021_g N_A_1728_125#_c_1849_n 8.62473e-19 $X=14.185 $Y=2.57
+ $X2=0 $Y2=0
cc_670 N_A_689_139#_c_598_n N_A_1728_125#_c_1808_n 0.0037442f $X=11.975 $Y=2.49
+ $X2=0 $Y2=0
cc_671 N_A_689_139#_c_575_n N_SET_B_M1027_g 0.00810283f $X=7.845 $Y=1.555 $X2=0
+ $Y2=0
cc_672 N_A_689_139#_M1025_g N_SET_B_c_2001_n 0.00737859f $X=8.205 $Y=0.945 $X2=0
+ $Y2=0
cc_673 N_A_689_139#_M1017_g N_SET_B_c_2001_n 0.00737859f $X=8.565 $Y=0.945 $X2=0
+ $Y2=0
cc_674 N_A_689_139#_M1021_g N_SET_B_M1043_g 0.0433479f $X=14.185 $Y=2.57 $X2=0
+ $Y2=0
cc_675 N_A_689_139#_c_600_n N_SET_B_M1043_g 0.015796f $X=14.04 $Y=2.095 $X2=0
+ $Y2=0
cc_676 N_A_689_139#_c_610_n N_SET_B_M1043_g 0.0040176f $X=13.27 $Y=2.095 $X2=0
+ $Y2=0
cc_677 N_A_689_139#_c_586_n N_SET_B_M1043_g 0.00170402f $X=14.205 $Y=1.745 $X2=0
+ $Y2=0
cc_678 N_A_689_139#_c_600_n N_SET_B_c_2005_n 9.58091e-19 $X=14.04 $Y=2.095 $X2=0
+ $Y2=0
cc_679 N_A_689_139#_c_587_n N_SET_B_c_2005_n 0.00966041f $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_680 N_A_689_139#_c_575_n N_SET_B_c_2008_n 0.00448628f $X=7.845 $Y=1.555 $X2=0
+ $Y2=0
cc_681 N_A_689_139#_c_600_n SET_B 0.0233962f $X=14.04 $Y=2.095 $X2=0 $Y2=0
cc_682 N_A_689_139#_c_586_n SET_B 0.0165476f $X=14.205 $Y=1.745 $X2=0 $Y2=0
cc_683 N_A_689_139#_c_587_n SET_B 3.28403e-19 $X=14.205 $Y=1.745 $X2=0 $Y2=0
cc_684 N_A_689_139#_M1021_g N_SET_B_c_2011_n 5.30612e-19 $X=14.185 $Y=2.57 $X2=0
+ $Y2=0
cc_685 N_A_689_139#_c_600_n N_SET_B_c_2011_n 0.00220015f $X=14.04 $Y=2.095 $X2=0
+ $Y2=0
cc_686 N_A_689_139#_c_586_n N_SET_B_c_2011_n 0.00160532f $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_687 N_A_689_139#_c_587_n N_SET_B_c_2011_n 0.020758f $X=14.205 $Y=1.745 $X2=0
+ $Y2=0
cc_688 N_A_689_139#_c_586_n CLK 0.00955767f $X=14.205 $Y=1.745 $X2=0 $Y2=0
cc_689 N_A_689_139#_c_576_n N_VPWR_c_2358_n 0.0310508f $X=7.93 $Y=2.905 $X2=0
+ $Y2=0
cc_690 N_A_689_139#_c_701_p N_VPWR_c_2358_n 0.0067793f $X=8.015 $Y=2.99 $X2=0
+ $Y2=0
cc_691 N_A_689_139#_M1005_g N_VPWR_c_2360_n 0.0054895f $X=5.155 $Y=2.885 $X2=0
+ $Y2=0
cc_692 N_A_689_139#_M1021_g N_VPWR_c_2365_n 0.00569155f $X=14.185 $Y=2.57 $X2=0
+ $Y2=0
cc_693 N_A_689_139#_c_647_p N_VPWR_c_2365_n 0.0402792f $X=8.525 $Y=2.99 $X2=0
+ $Y2=0
cc_694 N_A_689_139#_c_701_p N_VPWR_c_2365_n 0.0174653f $X=8.015 $Y=2.99 $X2=0
+ $Y2=0
cc_695 N_A_689_139#_M1005_g N_VPWR_c_2354_n 0.00672878f $X=5.155 $Y=2.885 $X2=0
+ $Y2=0
cc_696 N_A_689_139#_M1021_g N_VPWR_c_2354_n 0.00666363f $X=14.185 $Y=2.57 $X2=0
+ $Y2=0
cc_697 N_A_689_139#_c_647_p N_VPWR_c_2354_n 0.00557444f $X=8.525 $Y=2.99 $X2=0
+ $Y2=0
cc_698 N_A_689_139#_c_701_p N_VPWR_c_2354_n 0.0023256f $X=8.015 $Y=2.99 $X2=0
+ $Y2=0
cc_699 N_A_689_139#_M1010_d N_A_189_119#_c_2526_n 0.00483461f $X=3.575 $Y=1.795
+ $X2=0 $Y2=0
cc_700 N_A_689_139#_c_601_n N_A_189_119#_c_2526_n 0.0137542f $X=4.132 $Y=1.89
+ $X2=0 $Y2=0
cc_701 N_A_689_139#_c_602_n N_A_189_119#_c_2526_n 0.0274975f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_702 N_A_689_139#_c_603_n N_A_189_119#_c_2526_n 0.00167061f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_703 N_A_689_139#_M1010_d N_A_189_119#_c_2527_n 0.00131237f $X=3.575 $Y=1.795
+ $X2=0 $Y2=0
cc_704 N_A_689_139#_c_590_n N_A_189_119#_c_2528_n 0.00736363f $X=4.335 $Y=2.32
+ $X2=0 $Y2=0
cc_705 N_A_689_139#_c_601_n N_A_189_119#_c_2528_n 0.0120043f $X=4.132 $Y=1.89
+ $X2=0 $Y2=0
cc_706 N_A_689_139#_c_602_n N_A_189_119#_c_2528_n 0.00563374f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_707 N_A_689_139#_c_571_n N_A_189_119#_c_2520_n 0.0403191f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_708 N_A_689_139#_c_572_n N_A_189_119#_c_2520_n 0.00948186f $X=5.11 $Y=0.34
+ $X2=0 $Y2=0
cc_709 N_A_689_139#_c_579_n N_A_189_119#_c_2520_n 0.00273589f $X=4.015 $Y=0.42
+ $X2=0 $Y2=0
cc_710 N_A_689_139#_c_588_n N_A_189_119#_c_2520_n 4.004e-19 $X=3.85 $Y=0.18
+ $X2=0 $Y2=0
cc_711 N_A_689_139#_c_589_n N_A_189_119#_c_2521_n 0.00188541f $X=5.08 $Y=2.32
+ $X2=0 $Y2=0
cc_712 N_A_689_139#_c_602_n N_A_189_119#_c_2521_n 0.00221707f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_713 N_A_689_139#_c_603_n N_A_189_119#_c_2521_n 0.00196475f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_714 N_A_689_139#_c_571_n N_A_189_119#_c_2522_n 0.0120727f $X=3.585 $Y=0.905
+ $X2=0 $Y2=0
cc_715 N_A_689_139#_c_602_n N_A_189_119#_c_2522_n 0.0211864f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_716 N_A_689_139#_c_603_n N_A_189_119#_c_2522_n 0.0019752f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_717 N_A_689_139#_c_589_n N_A_189_119#_c_2523_n 0.0280016f $X=5.08 $Y=2.32
+ $X2=0 $Y2=0
cc_718 N_A_689_139#_M1005_g N_A_189_119#_c_2523_n 0.0120546f $X=5.155 $Y=2.885
+ $X2=0 $Y2=0
cc_719 N_A_689_139#_c_601_n N_A_189_119#_c_2523_n 0.02446f $X=4.132 $Y=1.89
+ $X2=0 $Y2=0
cc_720 N_A_689_139#_c_602_n N_A_189_119#_c_2523_n 0.02621f $X=4.17 $Y=1.89 $X2=0
+ $Y2=0
cc_721 N_A_689_139#_c_603_n N_A_189_119#_c_2523_n 0.0127461f $X=4.17 $Y=1.89
+ $X2=0 $Y2=0
cc_722 N_A_689_139#_c_576_n N_A_1541_125#_M1032_d 0.0187741f $X=7.93 $Y=2.905
+ $X2=0 $Y2=0
cc_723 N_A_689_139#_c_647_p N_A_1541_125#_M1032_d 0.0095041f $X=8.525 $Y=2.99
+ $X2=0 $Y2=0
cc_724 N_A_689_139#_c_701_p N_A_1541_125#_M1032_d 0.0062155f $X=8.015 $Y=2.99
+ $X2=0 $Y2=0
cc_725 N_A_689_139#_M1025_g N_A_1541_125#_c_2636_n 0.00742529f $X=8.205 $Y=0.945
+ $X2=0 $Y2=0
cc_726 N_A_689_139#_M1017_g N_A_1541_125#_c_2636_n 0.00127133f $X=8.565 $Y=0.945
+ $X2=0 $Y2=0
cc_727 N_A_689_139#_c_578_n N_A_1541_125#_c_2636_n 0.00698604f $X=8.695 $Y=0.68
+ $X2=0 $Y2=0
cc_728 N_A_689_139#_c_584_n N_A_1541_125#_c_2636_n 0.0121256f $X=8.64 $Y=1.41
+ $X2=0 $Y2=0
cc_729 N_A_689_139#_M1025_g N_A_1541_125#_c_2637_n 0.00423416f $X=8.205 $Y=0.945
+ $X2=0 $Y2=0
cc_730 N_A_689_139#_M1017_g N_A_1541_125#_c_2637_n 7.38556e-19 $X=8.565 $Y=0.945
+ $X2=0 $Y2=0
cc_731 N_A_689_139#_c_575_n N_A_1541_125#_c_2637_n 0.0137151f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_732 N_A_689_139#_c_576_n N_A_1541_125#_c_2637_n 0.0684096f $X=7.93 $Y=2.905
+ $X2=0 $Y2=0
cc_733 N_A_689_139#_c_647_p N_A_1541_125#_c_2637_n 0.00522009f $X=8.525 $Y=2.99
+ $X2=0 $Y2=0
cc_734 N_A_689_139#_c_583_n N_A_1541_125#_c_2637_n 0.0165541f $X=8.645 $Y=1.575
+ $X2=0 $Y2=0
cc_735 N_A_689_139#_c_584_n N_A_1541_125#_c_2637_n 0.0814284f $X=8.64 $Y=1.41
+ $X2=0 $Y2=0
cc_736 N_A_689_139#_M1025_g N_A_1541_125#_c_2653_n 0.00924903f $X=8.205 $Y=0.945
+ $X2=0 $Y2=0
cc_737 N_A_689_139#_M1017_g N_A_1541_125#_c_2653_n 9.65137e-19 $X=8.565 $Y=0.945
+ $X2=0 $Y2=0
cc_738 N_A_689_139#_c_575_n N_A_1541_125#_c_2653_n 0.0101338f $X=7.845 $Y=1.555
+ $X2=0 $Y2=0
cc_739 N_A_689_139#_c_584_n N_A_1541_125#_c_2653_n 0.0128807f $X=8.64 $Y=1.41
+ $X2=0 $Y2=0
cc_740 N_A_689_139#_c_647_p A_1712_451# 0.00229493f $X=8.525 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_741 N_A_689_139#_c_596_n A_1712_451# 0.00509309f $X=8.61 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_742 N_A_689_139#_c_724_p N_KAPWR_M1018_d 0.00743727f $X=13.185 $Y=2.31
+ $X2=-0.19 $Y2=-0.245
cc_743 N_A_689_139#_M1021_g N_KAPWR_c_2675_n 0.0130288f $X=14.185 $Y=2.57 $X2=0
+ $Y2=0
cc_744 N_A_689_139#_c_590_n N_KAPWR_c_2677_n 0.0010068f $X=4.335 $Y=2.32 $X2=0
+ $Y2=0
cc_745 N_A_689_139#_M1005_g N_KAPWR_c_2677_n 0.00685712f $X=5.155 $Y=2.885 $X2=0
+ $Y2=0
cc_746 N_A_689_139#_M1021_g N_KAPWR_c_2677_n 0.00463752f $X=14.185 $Y=2.57 $X2=0
+ $Y2=0
cc_747 N_A_689_139#_c_576_n N_KAPWR_c_2677_n 0.0219785f $X=7.93 $Y=2.905 $X2=0
+ $Y2=0
cc_748 N_A_689_139#_c_647_p N_KAPWR_c_2677_n 0.0195076f $X=8.525 $Y=2.99 $X2=0
+ $Y2=0
cc_749 N_A_689_139#_c_701_p N_KAPWR_c_2677_n 0.00615246f $X=8.015 $Y=2.99 $X2=0
+ $Y2=0
cc_750 N_A_689_139#_c_596_n N_KAPWR_c_2677_n 0.020636f $X=8.61 $Y=2.905 $X2=0
+ $Y2=0
cc_751 N_A_689_139#_c_598_n N_KAPWR_c_2677_n 0.0754478f $X=11.975 $Y=2.49 $X2=0
+ $Y2=0
cc_752 N_A_689_139#_c_599_n N_KAPWR_c_2677_n 0.00537759f $X=9.485 $Y=2.49 $X2=0
+ $Y2=0
cc_753 N_A_689_139#_c_724_p N_KAPWR_c_2677_n 0.00944884f $X=13.185 $Y=2.31 $X2=0
+ $Y2=0
cc_754 N_A_689_139#_c_600_n N_KAPWR_c_2677_n 0.00326147f $X=14.04 $Y=2.095 $X2=0
+ $Y2=0
cc_755 N_A_689_139#_c_601_n N_KAPWR_c_2677_n 0.00170269f $X=4.132 $Y=1.89 $X2=0
+ $Y2=0
cc_756 N_A_689_139#_c_725_p N_KAPWR_c_2677_n 0.00522441f $X=12.06 $Y=2.31 $X2=0
+ $Y2=0
cc_757 N_A_689_139#_c_610_n N_KAPWR_c_2677_n 9.86236e-19 $X=13.27 $Y=2.095 $X2=0
+ $Y2=0
cc_758 N_A_689_139#_c_586_n N_KAPWR_c_2677_n 5.25934e-19 $X=14.205 $Y=1.745
+ $X2=0 $Y2=0
cc_759 N_A_689_139#_c_600_n A_2658_414# 0.00203746f $X=14.04 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_760 N_A_689_139#_c_610_n A_2658_414# 0.00288915f $X=13.27 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_761 N_A_689_139#_c_571_n N_VGND_c_2835_n 0.020482f $X=3.585 $Y=0.905 $X2=0
+ $Y2=0
cc_762 N_A_689_139#_c_579_n N_VGND_c_2835_n 0.0287821f $X=4.015 $Y=0.42 $X2=0
+ $Y2=0
cc_763 N_A_689_139#_c_588_n N_VGND_c_2835_n 0.00437546f $X=3.85 $Y=0.18 $X2=0
+ $Y2=0
cc_764 N_A_689_139#_c_567_n N_VGND_c_2836_n 0.00107184f $X=4.83 $Y=0.18 $X2=0
+ $Y2=0
cc_765 N_A_689_139#_c_572_n N_VGND_c_2836_n 0.0131487f $X=5.11 $Y=0.34 $X2=0
+ $Y2=0
cc_766 N_A_689_139#_c_573_n N_VGND_c_2836_n 0.00549917f $X=5.195 $Y=1.545 $X2=0
+ $Y2=0
cc_767 N_A_689_139#_c_572_n N_VGND_c_2850_n 0.0119531f $X=5.11 $Y=0.34 $X2=0
+ $Y2=0
cc_768 N_A_689_139#_c_579_n N_VGND_c_2850_n 0.109123f $X=4.015 $Y=0.42 $X2=0
+ $Y2=0
cc_769 N_A_689_139#_c_588_n N_VGND_c_2850_n 0.0281467f $X=3.85 $Y=0.18 $X2=0
+ $Y2=0
cc_770 N_A_689_139#_c_567_n N_VGND_c_2854_n 0.0240041f $X=4.83 $Y=0.18 $X2=0
+ $Y2=0
cc_771 N_A_689_139#_c_572_n N_VGND_c_2854_n 0.00660921f $X=5.11 $Y=0.34 $X2=0
+ $Y2=0
cc_772 N_A_689_139#_c_579_n N_VGND_c_2854_n 0.0583693f $X=4.015 $Y=0.42 $X2=0
+ $Y2=0
cc_773 N_A_689_139#_c_588_n N_VGND_c_2854_n 0.0101308f $X=3.85 $Y=0.18 $X2=0
+ $Y2=0
cc_774 N_A_689_139#_c_572_n A_996_73# 0.00720528f $X=5.11 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_775 N_A_689_139#_c_573_n A_996_73# 0.00837648f $X=5.195 $Y=1.545 $X2=-0.19
+ $Y2=-0.245
cc_776 N_A_659_113#_c_908_n N_A_1068_21#_c_1248_n 0.00378015f $X=5.78 $Y=0.76
+ $X2=0 $Y2=0
cc_777 N_A_659_113#_c_909_n N_A_1068_21#_c_1248_n 0.00310765f $X=6.05 $Y=0.675
+ $X2=0 $Y2=0
cc_778 N_A_659_113#_c_905_n N_A_1068_21#_c_1249_n 0.00593849f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_779 N_A_659_113#_c_907_n N_A_1068_21#_c_1249_n 0.0119934f $X=5.965 $Y=0.76
+ $X2=0 $Y2=0
cc_780 N_A_659_113#_c_908_n N_A_1068_21#_c_1249_n 0.00680324f $X=5.78 $Y=0.76
+ $X2=0 $Y2=0
cc_781 N_A_659_113#_c_901_n N_A_1068_21#_c_1250_n 0.00524977f $X=5.45 $Y=1.3
+ $X2=0 $Y2=0
cc_782 N_A_659_113#_c_905_n N_A_1068_21#_c_1250_n 0.00114094f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_783 N_A_659_113#_c_906_n N_A_1068_21#_c_1250_n 0.0213685f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_784 N_A_659_113#_c_908_n N_A_1068_21#_c_1250_n 9.11332e-19 $X=5.78 $Y=0.76
+ $X2=0 $Y2=0
cc_785 N_A_659_113#_c_905_n N_A_1068_21#_c_1251_n 0.00362021f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_786 N_A_659_113#_c_906_n N_A_1068_21#_c_1251_n 0.014552f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_787 N_A_659_113#_c_907_n N_A_1068_21#_c_1251_n 0.00682375f $X=5.965 $Y=0.76
+ $X2=0 $Y2=0
cc_788 N_A_659_113#_c_910_n N_A_1068_21#_c_1251_n 0.00306779f $X=6.725 $Y=0.34
+ $X2=0 $Y2=0
cc_789 N_A_659_113#_c_905_n N_A_1068_21#_c_1252_n 0.0192372f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_790 N_A_659_113#_c_906_n N_A_1068_21#_c_1252_n 6.46553e-19 $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_791 N_A_659_113#_c_907_n N_A_1068_21#_c_1252_n 0.0113227f $X=5.965 $Y=0.76
+ $X2=0 $Y2=0
cc_792 N_A_659_113#_c_910_n N_A_1068_21#_c_1252_n 0.00489653f $X=6.725 $Y=0.34
+ $X2=0 $Y2=0
cc_793 N_A_659_113#_c_912_n N_A_1068_21#_c_1252_n 0.00901783f $X=6.81 $Y=1.13
+ $X2=0 $Y2=0
cc_794 N_A_659_113#_c_914_n N_A_1068_21#_c_1252_n 0.0149552f $X=6.895 $Y=1.215
+ $X2=0 $Y2=0
cc_795 N_A_659_113#_c_905_n N_A_1068_21#_c_1253_n 0.00589307f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_796 N_A_659_113#_c_907_n N_A_1068_21#_c_1253_n 0.0141465f $X=5.965 $Y=0.76
+ $X2=0 $Y2=0
cc_797 N_A_659_113#_c_909_n N_A_1068_21#_c_1253_n 0.00605232f $X=6.05 $Y=0.675
+ $X2=0 $Y2=0
cc_798 N_A_659_113#_c_910_n N_A_1068_21#_c_1253_n 0.0168013f $X=6.725 $Y=0.34
+ $X2=0 $Y2=0
cc_799 N_A_659_113#_c_912_n N_A_1068_21#_c_1253_n 0.019168f $X=6.81 $Y=1.13
+ $X2=0 $Y2=0
cc_800 N_A_659_113#_M1034_g N_A_1068_21#_c_1257_n 0.0569159f $X=5.585 $Y=2.885
+ $X2=0 $Y2=0
cc_801 N_A_659_113#_M1034_g N_A_1068_21#_c_1258_n 8.23572e-19 $X=5.585 $Y=2.885
+ $X2=0 $Y2=0
cc_802 N_A_659_113#_M1034_g N_A_1068_21#_c_1254_n 0.0210267f $X=5.585 $Y=2.885
+ $X2=0 $Y2=0
cc_803 N_A_659_113#_c_906_n N_A_1068_21#_c_1254_n 0.00547445f $X=5.615 $Y=1.29
+ $X2=0 $Y2=0
cc_804 N_A_659_113#_c_909_n N_A_887_139#_M1038_g 0.00259659f $X=6.05 $Y=0.675
+ $X2=0 $Y2=0
cc_805 N_A_659_113#_c_910_n N_A_887_139#_M1038_g 0.0114507f $X=6.725 $Y=0.34
+ $X2=0 $Y2=0
cc_806 N_A_659_113#_c_912_n N_A_887_139#_M1038_g 0.00379658f $X=6.81 $Y=1.13
+ $X2=0 $Y2=0
cc_807 N_A_659_113#_c_914_n N_A_887_139#_M1038_g 0.0013169f $X=6.895 $Y=1.215
+ $X2=0 $Y2=0
cc_808 N_A_659_113#_c_913_n N_A_887_139#_M1040_g 0.00766355f $X=7.535 $Y=1.215
+ $X2=0 $Y2=0
cc_809 N_A_659_113#_c_915_n N_A_887_139#_M1040_g 0.0189616f $X=7.62 $Y=1.13
+ $X2=0 $Y2=0
cc_810 N_A_659_113#_c_930_n N_A_887_139#_M1032_g 0.00587112f $X=8.485 $Y=2.145
+ $X2=0 $Y2=0
cc_811 N_A_659_113#_c_900_n N_A_887_139#_c_1345_n 0.00166369f $X=4.36 $Y=1.225
+ $X2=0 $Y2=0
cc_812 N_A_659_113#_c_901_n N_A_887_139#_c_1345_n 0.0139479f $X=5.45 $Y=1.3
+ $X2=0 $Y2=0
cc_813 N_A_659_113#_M1034_g N_A_887_139#_c_1345_n 0.00492127f $X=5.585 $Y=2.885
+ $X2=0 $Y2=0
cc_814 N_A_659_113#_c_901_n N_A_887_139#_c_1352_n 0.00431959f $X=5.45 $Y=1.3
+ $X2=0 $Y2=0
cc_815 N_A_659_113#_M1034_g N_A_887_139#_c_1354_n 0.0243953f $X=5.585 $Y=2.885
+ $X2=0 $Y2=0
cc_816 N_A_659_113#_c_932_n N_A_887_139#_c_1346_n 0.00587112f $X=8.56 $Y=2.07
+ $X2=0 $Y2=0
cc_817 N_A_659_113#_c_913_n N_A_887_139#_c_1346_n 0.00106408f $X=7.535 $Y=1.215
+ $X2=0 $Y2=0
cc_818 N_A_659_113#_c_900_n N_A_887_139#_c_1347_n 0.00775612f $X=4.36 $Y=1.225
+ $X2=0 $Y2=0
cc_819 N_A_659_113#_c_901_n N_A_887_139#_c_1347_n 0.0115924f $X=5.45 $Y=1.3
+ $X2=0 $Y2=0
cc_820 N_A_659_113#_c_901_n N_A_887_139#_c_1359_n 6.02688e-19 $X=5.45 $Y=1.3
+ $X2=0 $Y2=0
cc_821 N_A_659_113#_M1034_g N_A_887_139#_c_1359_n 0.00487959f $X=5.585 $Y=2.885
+ $X2=0 $Y2=0
cc_822 N_A_659_113#_M1034_g N_A_887_139#_c_1360_n 0.00941048f $X=5.585 $Y=2.885
+ $X2=0 $Y2=0
cc_823 N_A_659_113#_c_921_n N_A_1972_99#_M1041_d 0.0117064f $X=13.185 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_824 N_A_659_113#_M1050_g N_A_1972_99#_M1046_g 0.063683f $X=9.575 $Y=0.835
+ $X2=0 $Y2=0
cc_825 N_A_659_113#_c_916_n N_A_1972_99#_M1046_g 0.00366331f $X=10.085 $Y=0.34
+ $X2=0 $Y2=0
cc_826 N_A_659_113#_c_918_n N_A_1972_99#_M1046_g 0.010889f $X=10.17 $Y=1.545
+ $X2=0 $Y2=0
cc_827 N_A_659_113#_c_918_n N_A_1972_99#_c_1474_n 0.00431555f $X=10.17 $Y=1.545
+ $X2=0 $Y2=0
cc_828 N_A_659_113#_c_940_n N_A_1972_99#_c_1474_n 0.0179191f $X=10.25 $Y=1.98
+ $X2=0 $Y2=0
cc_829 N_A_659_113#_c_926_n N_A_1972_99#_c_1474_n 0.00196658f $X=10.25 $Y=1.63
+ $X2=0 $Y2=0
cc_830 N_A_659_113#_c_936_n N_A_1972_99#_c_1475_n 0.00893448f $X=10.085 $Y=2.07
+ $X2=0 $Y2=0
cc_831 N_A_659_113#_c_918_n N_A_1972_99#_M1006_g 0.0177273f $X=10.17 $Y=1.545
+ $X2=0 $Y2=0
cc_832 N_A_659_113#_c_919_n N_A_1972_99#_c_1477_n 0.00924942f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_833 N_A_659_113#_c_926_n N_A_1972_99#_c_1477_n 0.0024683f $X=10.25 $Y=1.63
+ $X2=0 $Y2=0
cc_834 N_A_659_113#_c_918_n N_A_1972_99#_c_1478_n 0.0053946f $X=10.17 $Y=1.545
+ $X2=0 $Y2=0
cc_835 N_A_659_113#_c_926_n N_A_1972_99#_c_1478_n 0.00787378f $X=10.25 $Y=1.63
+ $X2=0 $Y2=0
cc_836 N_A_659_113#_c_919_n N_A_1972_99#_c_1488_n 0.0359166f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_837 N_A_659_113#_c_919_n N_A_1972_99#_c_1489_n 0.0624386f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_838 N_A_659_113#_c_920_n N_A_1972_99#_c_1531_n 0.0213763f $X=12.59 $Y=1.545
+ $X2=0 $Y2=0
cc_839 N_A_659_113#_c_921_n N_A_1972_99#_c_1531_n 0.0136682f $X=13.185 $Y=0.68
+ $X2=0 $Y2=0
cc_840 N_A_659_113#_c_927_n N_A_1972_99#_c_1531_n 0.00998544f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_841 N_A_659_113#_c_919_n N_A_1972_99#_c_1480_n 0.0135857f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_842 N_A_659_113#_c_920_n N_A_1972_99#_c_1480_n 0.00958428f $X=12.59 $Y=1.545
+ $X2=0 $Y2=0
cc_843 N_A_659_113#_c_921_n N_A_1972_99#_c_1481_n 0.0059505f $X=13.185 $Y=0.68
+ $X2=0 $Y2=0
cc_844 N_A_659_113#_c_922_n N_A_1972_99#_c_1481_n 0.0524304f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_845 N_A_659_113#_c_923_n N_A_1972_99#_c_1481_n 0.00736571f $X=15.405 $Y=0.72
+ $X2=0 $Y2=0
cc_846 N_A_659_113#_c_924_n N_A_1972_99#_c_1481_n 0.0127363f $X=14.255 $Y=0.72
+ $X2=0 $Y2=0
cc_847 N_A_659_113#_c_927_n N_A_1972_99#_c_1481_n 0.012997f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_848 N_A_659_113#_c_939_n N_A_1972_99#_c_1491_n 0.0145039f $X=10.25 $Y=1.98
+ $X2=0 $Y2=0
cc_849 N_A_659_113#_c_940_n N_A_1972_99#_c_1491_n 0.00104596f $X=10.25 $Y=1.98
+ $X2=0 $Y2=0
cc_850 N_A_659_113#_c_919_n N_A_1972_99#_c_1491_n 0.0242156f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_851 N_A_659_113#_c_919_n N_A_1972_99#_c_1492_n 0.00126186f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_852 N_A_659_113#_c_919_n N_A_1972_99#_c_1493_n 0.0248805f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_853 N_A_659_113#_c_920_n N_A_1972_99#_c_1482_n 0.0137075f $X=12.59 $Y=1.545
+ $X2=0 $Y2=0
cc_854 N_A_659_113#_c_923_n N_A_1972_99#_c_1483_n 0.0232047f $X=15.405 $Y=0.72
+ $X2=0 $Y2=0
cc_855 N_A_659_113#_c_924_n N_A_1972_99#_c_1483_n 0.0022547f $X=14.255 $Y=0.72
+ $X2=0 $Y2=0
cc_856 N_A_659_113#_c_925_n N_A_1972_99#_c_1483_n 0.00374734f $X=15.49 $Y=1.9
+ $X2=0 $Y2=0
cc_857 N_A_659_113#_c_923_n N_A_1972_99#_c_1484_n 0.00230176f $X=15.405 $Y=0.72
+ $X2=0 $Y2=0
cc_858 N_A_659_113#_c_939_n N_A_1972_99#_c_1485_n 0.00471888f $X=10.25 $Y=1.98
+ $X2=0 $Y2=0
cc_859 N_A_659_113#_c_940_n N_A_1972_99#_c_1485_n 0.0178339f $X=10.25 $Y=1.98
+ $X2=0 $Y2=0
cc_860 N_A_659_113#_c_919_n N_A_1972_99#_c_1485_n 0.0104909f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_861 N_A_659_113#_c_919_n N_A_2216_99#_c_1617_n 0.00154805f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_862 N_A_659_113#_c_921_n N_A_2216_99#_c_1618_n 0.00143288f $X=13.185 $Y=0.68
+ $X2=0 $Y2=0
cc_863 N_A_659_113#_c_927_n N_A_2216_99#_c_1618_n 0.00347622f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_864 N_A_659_113#_c_922_n N_A_2216_99#_c_1620_n 0.00947797f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_865 N_A_659_113#_c_924_n N_A_2216_99#_c_1620_n 6.0417e-19 $X=14.255 $Y=0.72
+ $X2=0 $Y2=0
cc_866 N_A_659_113#_c_927_n N_A_2216_99#_c_1620_n 0.00945665f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_867 N_A_659_113#_c_919_n N_A_2216_99#_c_1621_n 0.0535722f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_868 N_A_659_113#_c_920_n N_A_2216_99#_c_1621_n 0.0211825f $X=12.59 $Y=1.545
+ $X2=0 $Y2=0
cc_869 N_A_659_113#_c_919_n N_A_2216_99#_c_1622_n 0.00244803f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_870 N_A_659_113#_c_920_n N_A_2216_99#_c_1623_n 0.00816707f $X=12.59 $Y=1.545
+ $X2=0 $Y2=0
cc_871 N_A_659_113#_c_921_n N_A_2216_99#_c_1624_n 0.0338531f $X=13.185 $Y=0.68
+ $X2=0 $Y2=0
cc_872 N_A_659_113#_c_1112_p N_A_2216_99#_c_1624_n 0.0120034f $X=12.675 $Y=0.68
+ $X2=0 $Y2=0
cc_873 N_A_659_113#_c_922_n N_A_2216_99#_c_1624_n 0.0058169f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_874 N_A_659_113#_c_927_n N_A_2216_99#_c_1624_n 0.0127788f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_875 N_A_659_113#_M1015_s N_A_2216_99#_c_1626_n 0.00441335f $X=14.73 $Y=0.36
+ $X2=0 $Y2=0
cc_876 N_A_659_113#_c_922_n N_A_2216_99#_c_1626_n 0.0083594f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_877 N_A_659_113#_c_923_n N_A_2216_99#_c_1626_n 0.0816243f $X=15.405 $Y=0.72
+ $X2=0 $Y2=0
cc_878 N_A_659_113#_c_924_n N_A_2216_99#_c_1626_n 0.0119335f $X=14.255 $Y=0.72
+ $X2=0 $Y2=0
cc_879 N_A_659_113#_c_923_n N_A_2216_99#_c_1627_n 0.0197346f $X=15.405 $Y=0.72
+ $X2=0 $Y2=0
cc_880 N_A_659_113#_c_925_n N_A_2216_99#_c_1627_n 0.00243153f $X=15.49 $Y=1.9
+ $X2=0 $Y2=0
cc_881 N_A_659_113#_c_925_n N_A_2216_99#_c_1629_n 0.0132531f $X=15.49 $Y=1.9
+ $X2=0 $Y2=0
cc_882 N_A_659_113#_c_922_n N_A_2216_99#_c_1632_n 0.0254762f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_883 N_A_659_113#_c_924_n N_A_2216_99#_c_1632_n 0.00757151f $X=14.255 $Y=0.72
+ $X2=0 $Y2=0
cc_884 N_A_659_113#_c_927_n N_A_2216_99#_c_1632_n 0.00964069f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_885 N_A_659_113#_c_921_n N_A_2216_99#_c_1633_n 3.81406e-19 $X=13.185 $Y=0.68
+ $X2=0 $Y2=0
cc_886 N_A_659_113#_c_922_n N_A_2216_99#_c_1633_n 0.00682232f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_887 N_A_659_113#_c_924_n N_A_2216_99#_c_1633_n 9.67451e-19 $X=14.255 $Y=0.72
+ $X2=0 $Y2=0
cc_888 N_A_659_113#_c_927_n N_A_2216_99#_c_1633_n 0.00805219f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_889 N_A_659_113#_c_919_n N_A_2216_99#_c_1634_n 0.00346708f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_890 N_A_659_113#_c_919_n N_A_1728_125#_c_1793_n 0.0116721f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_891 N_A_659_113#_c_919_n N_A_1728_125#_M1051_g 0.012025f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_892 N_A_659_113#_c_920_n N_A_1728_125#_M1051_g 0.00446821f $X=12.59 $Y=1.545
+ $X2=0 $Y2=0
cc_893 N_A_659_113#_c_919_n N_A_1728_125#_M1041_g 0.00612585f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_894 N_A_659_113#_c_920_n N_A_1728_125#_M1041_g 0.017158f $X=12.59 $Y=1.545
+ $X2=0 $Y2=0
cc_895 N_A_659_113#_c_1112_p N_A_1728_125#_M1041_g 0.00703537f $X=12.675 $Y=0.68
+ $X2=0 $Y2=0
cc_896 N_A_659_113#_c_927_n N_A_1728_125#_M1041_g 0.00145659f $X=13.27 $Y=0.68
+ $X2=0 $Y2=0
cc_897 N_A_659_113#_c_919_n N_A_1728_125#_c_1799_n 9.32779e-19 $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_898 N_A_659_113#_c_930_n N_A_1728_125#_c_1800_n 3.17938e-19 $X=8.485 $Y=2.145
+ $X2=0 $Y2=0
cc_899 N_A_659_113#_c_933_n N_A_1728_125#_c_1800_n 0.0027653f $X=8.845 $Y=2.145
+ $X2=0 $Y2=0
cc_900 N_A_659_113#_c_934_n N_A_1728_125#_c_1800_n 0.00239323f $X=9.5 $Y=2.07
+ $X2=0 $Y2=0
cc_901 N_A_659_113#_c_933_n N_A_1728_125#_c_1823_n 0.0031862f $X=8.845 $Y=2.145
+ $X2=0 $Y2=0
cc_902 N_A_659_113#_c_933_n N_A_1728_125#_c_1825_n 0.00320175f $X=8.845 $Y=2.145
+ $X2=0 $Y2=0
cc_903 N_A_659_113#_c_934_n N_A_1728_125#_c_1801_n 0.00390018f $X=9.5 $Y=2.07
+ $X2=0 $Y2=0
cc_904 N_A_659_113#_M1039_d N_A_1728_125#_c_1802_n 0.00395257f $X=15.46 $Y=1.92
+ $X2=0 $Y2=0
cc_905 N_A_659_113#_c_944_n N_A_1728_125#_c_1802_n 0.0173041f $X=15.6 $Y=2.065
+ $X2=0 $Y2=0
cc_906 N_A_659_113#_M1050_g N_A_1728_125#_c_1833_n 0.00155347f $X=9.575 $Y=0.835
+ $X2=0 $Y2=0
cc_907 N_A_659_113#_c_933_n N_A_1728_125#_c_1788_n 0.00216306f $X=8.845 $Y=2.145
+ $X2=0 $Y2=0
cc_908 N_A_659_113#_c_934_n N_A_1728_125#_c_1788_n 0.0152177f $X=9.5 $Y=2.07
+ $X2=0 $Y2=0
cc_909 N_A_659_113#_M1050_g N_A_1728_125#_c_1788_n 0.00317421f $X=9.575 $Y=0.835
+ $X2=0 $Y2=0
cc_910 N_A_659_113#_c_910_n N_SET_B_M1003_g 0.00310286f $X=6.725 $Y=0.34 $X2=0
+ $Y2=0
cc_911 N_A_659_113#_c_912_n N_SET_B_M1003_g 0.00470401f $X=6.81 $Y=1.13 $X2=0
+ $Y2=0
cc_912 N_A_659_113#_c_913_n N_SET_B_M1003_g 0.0152388f $X=7.535 $Y=1.215 $X2=0
+ $Y2=0
cc_913 N_A_659_113#_c_915_n N_SET_B_M1003_g 7.92541e-19 $X=7.62 $Y=1.13 $X2=0
+ $Y2=0
cc_914 N_A_659_113#_M1050_g N_SET_B_c_2001_n 0.00737859f $X=9.575 $Y=0.835 $X2=0
+ $Y2=0
cc_915 N_A_659_113#_c_916_n N_SET_B_c_2001_n 0.0497796f $X=10.085 $Y=0.34 $X2=0
+ $Y2=0
cc_916 N_A_659_113#_c_917_n N_SET_B_c_2001_n 0.00176618f $X=7.705 $Y=0.34 $X2=0
+ $Y2=0
cc_917 N_A_659_113#_c_916_n N_SET_B_M1008_g 0.00317758f $X=10.085 $Y=0.34 $X2=0
+ $Y2=0
cc_918 N_A_659_113#_c_918_n N_SET_B_M1008_g 0.00170032f $X=10.17 $Y=1.545 $X2=0
+ $Y2=0
cc_919 N_A_659_113#_c_922_n N_SET_B_c_2004_n 2.89005e-19 $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_920 N_A_659_113#_c_922_n N_SET_B_c_2006_n 0.00584839f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_921 N_A_659_113#_c_922_n N_SET_B_c_2007_n 0.00481619f $X=14.085 $Y=0.985
+ $X2=0 $Y2=0
cc_922 N_A_659_113#_c_923_n N_SET_B_c_2007_n 0.00260961f $X=15.405 $Y=0.72 $X2=0
+ $Y2=0
cc_923 N_A_659_113#_c_924_n N_SET_B_c_2007_n 0.019941f $X=14.255 $Y=0.72 $X2=0
+ $Y2=0
cc_924 N_A_659_113#_c_913_n N_SET_B_c_2008_n 0.00184328f $X=7.535 $Y=1.215 $X2=0
+ $Y2=0
cc_925 N_A_659_113#_c_923_n N_CLK_M1015_g 0.0182779f $X=15.405 $Y=0.72 $X2=0
+ $Y2=0
cc_926 N_A_659_113#_c_925_n N_CLK_M1015_g 0.00697695f $X=15.49 $Y=1.9 $X2=0
+ $Y2=0
cc_927 N_A_659_113#_c_925_n N_CLK_M1039_g 0.00443976f $X=15.49 $Y=1.9 $X2=0
+ $Y2=0
cc_928 N_A_659_113#_c_944_n N_CLK_M1039_g 0.00420665f $X=15.6 $Y=2.065 $X2=0
+ $Y2=0
cc_929 N_A_659_113#_c_923_n CLK 0.0135924f $X=15.405 $Y=0.72 $X2=0 $Y2=0
cc_930 N_A_659_113#_c_925_n CLK 0.0520405f $X=15.49 $Y=1.9 $X2=0 $Y2=0
cc_931 N_A_659_113#_c_944_n CLK 0.0192048f $X=15.6 $Y=2.065 $X2=0 $Y2=0
cc_932 N_A_659_113#_c_923_n N_CLK_c_2123_n 0.00448813f $X=15.405 $Y=0.72 $X2=0
+ $Y2=0
cc_933 N_A_659_113#_c_925_n N_CLK_c_2123_n 0.00921243f $X=15.49 $Y=1.9 $X2=0
+ $Y2=0
cc_934 N_A_659_113#_c_923_n N_SLEEP_B_M1014_g 0.00636876f $X=15.405 $Y=0.72
+ $X2=0 $Y2=0
cc_935 N_A_659_113#_c_925_n N_SLEEP_B_M1014_g 0.00189512f $X=15.49 $Y=1.9 $X2=0
+ $Y2=0
cc_936 N_A_659_113#_c_925_n N_SLEEP_B_M1026_g 0.00269524f $X=15.49 $Y=1.9 $X2=0
+ $Y2=0
cc_937 N_A_659_113#_c_944_n N_SLEEP_B_M1026_g 0.00425981f $X=15.6 $Y=2.065 $X2=0
+ $Y2=0
cc_938 N_A_659_113#_c_923_n N_SLEEP_B_M1049_g 2.08867e-19 $X=15.405 $Y=0.72
+ $X2=0 $Y2=0
cc_939 N_A_659_113#_c_925_n N_SLEEP_B_c_2168_n 0.0305677f $X=15.49 $Y=1.9 $X2=0
+ $Y2=0
cc_940 N_A_659_113#_c_944_n N_SLEEP_B_c_2168_n 0.0102334f $X=15.6 $Y=2.065 $X2=0
+ $Y2=0
cc_941 N_A_659_113#_c_925_n N_SLEEP_B_c_2169_n 0.0129652f $X=15.49 $Y=1.9 $X2=0
+ $Y2=0
cc_942 N_A_659_113#_c_944_n N_SLEEP_B_c_2169_n 0.00249232f $X=15.6 $Y=2.065
+ $X2=0 $Y2=0
cc_943 N_A_659_113#_c_897_n N_VPWR_c_2356_n 0.00787879f $X=3.5 $Y=1.375 $X2=0
+ $Y2=0
cc_944 N_A_659_113#_M1034_g N_VPWR_c_2357_n 0.0024931f $X=5.585 $Y=2.885 $X2=0
+ $Y2=0
cc_945 N_A_659_113#_c_897_n N_VPWR_c_2360_n 0.00345047f $X=3.5 $Y=1.375 $X2=0
+ $Y2=0
cc_946 N_A_659_113#_M1034_g N_VPWR_c_2360_n 0.0054895f $X=5.585 $Y=2.885 $X2=0
+ $Y2=0
cc_947 N_A_659_113#_c_930_n N_VPWR_c_2365_n 0.00357828f $X=8.485 $Y=2.145 $X2=0
+ $Y2=0
cc_948 N_A_659_113#_c_933_n N_VPWR_c_2365_n 0.00557384f $X=8.845 $Y=2.145 $X2=0
+ $Y2=0
cc_949 N_A_659_113#_c_897_n N_VPWR_c_2354_n 8.74848e-19 $X=3.5 $Y=1.375 $X2=0
+ $Y2=0
cc_950 N_A_659_113#_M1034_g N_VPWR_c_2354_n 0.00524789f $X=5.585 $Y=2.885 $X2=0
+ $Y2=0
cc_951 N_A_659_113#_c_930_n N_VPWR_c_2354_n 0.00541146f $X=8.485 $Y=2.145 $X2=0
+ $Y2=0
cc_952 N_A_659_113#_c_933_n N_VPWR_c_2354_n 0.00651507f $X=8.845 $Y=2.145 $X2=0
+ $Y2=0
cc_953 N_A_659_113#_c_897_n N_A_189_119#_c_2526_n 0.0122567f $X=3.5 $Y=1.375
+ $X2=0 $Y2=0
cc_954 N_A_659_113#_c_897_n N_A_189_119#_c_2527_n 0.0084934f $X=3.5 $Y=1.375
+ $X2=0 $Y2=0
cc_955 N_A_659_113#_c_897_n N_A_189_119#_c_2529_n 0.00369912f $X=3.5 $Y=1.375
+ $X2=0 $Y2=0
cc_956 N_A_659_113#_c_896_n N_A_189_119#_c_2520_n 0.0010368f $X=3.37 $Y=1.225
+ $X2=0 $Y2=0
cc_957 N_A_659_113#_c_898_n N_A_189_119#_c_2520_n 0.0171092f $X=4.285 $Y=1.3
+ $X2=0 $Y2=0
cc_958 N_A_659_113#_c_900_n N_A_189_119#_c_2520_n 0.00290404f $X=4.36 $Y=1.225
+ $X2=0 $Y2=0
cc_959 N_A_659_113#_c_898_n N_A_189_119#_c_2521_n 0.00734883f $X=4.285 $Y=1.3
+ $X2=0 $Y2=0
cc_960 N_A_659_113#_c_904_n N_A_189_119#_c_2521_n 0.00447261f $X=4.36 $Y=1.3
+ $X2=0 $Y2=0
cc_961 N_A_659_113#_c_897_n N_A_189_119#_c_2522_n 8.97762e-19 $X=3.5 $Y=1.375
+ $X2=0 $Y2=0
cc_962 N_A_659_113#_c_915_n N_A_1541_125#_c_2636_n 0.0364485f $X=7.62 $Y=1.13
+ $X2=0 $Y2=0
cc_963 N_A_659_113#_c_916_n N_A_1541_125#_c_2636_n 0.0206202f $X=10.085 $Y=0.34
+ $X2=0 $Y2=0
cc_964 N_A_659_113#_c_932_n N_A_1541_125#_c_2637_n 0.00359868f $X=8.56 $Y=2.07
+ $X2=0 $Y2=0
cc_965 N_A_659_113#_c_913_n N_A_1541_125#_c_2637_n 0.00114274f $X=7.535 $Y=1.215
+ $X2=0 $Y2=0
cc_966 N_A_659_113#_c_913_n N_A_1541_125#_c_2653_n 0.0114081f $X=7.535 $Y=1.215
+ $X2=0 $Y2=0
cc_967 N_A_659_113#_c_915_n N_A_1541_125#_c_2653_n 0.00257278f $X=7.62 $Y=1.13
+ $X2=0 $Y2=0
cc_968 N_A_659_113#_c_916_n N_A_1541_125#_c_2653_n 0.00471805f $X=10.085 $Y=0.34
+ $X2=0 $Y2=0
cc_969 N_A_659_113#_c_897_n N_KAPWR_c_2677_n 0.0124692f $X=3.5 $Y=1.375 $X2=0
+ $Y2=0
cc_970 N_A_659_113#_M1034_g N_KAPWR_c_2677_n 0.00452376f $X=5.585 $Y=2.885 $X2=0
+ $Y2=0
cc_971 N_A_659_113#_c_930_n N_KAPWR_c_2677_n 0.00787153f $X=8.485 $Y=2.145 $X2=0
+ $Y2=0
cc_972 N_A_659_113#_c_933_n N_KAPWR_c_2677_n 0.00779525f $X=8.845 $Y=2.145 $X2=0
+ $Y2=0
cc_973 N_A_659_113#_c_934_n N_KAPWR_c_2677_n 0.0032954f $X=9.5 $Y=2.07 $X2=0
+ $Y2=0
cc_974 N_A_659_113#_c_913_n N_VGND_M1003_d 0.00827774f $X=7.535 $Y=1.215 $X2=0
+ $Y2=0
cc_975 N_A_659_113#_c_896_n N_VGND_c_2835_n 0.00276581f $X=3.37 $Y=1.225 $X2=0
+ $Y2=0
cc_976 N_A_659_113#_c_907_n N_VGND_c_2836_n 0.00108678f $X=5.965 $Y=0.76 $X2=0
+ $Y2=0
cc_977 N_A_659_113#_c_908_n N_VGND_c_2836_n 0.0246151f $X=5.78 $Y=0.76 $X2=0
+ $Y2=0
cc_978 N_A_659_113#_c_909_n N_VGND_c_2836_n 0.00630512f $X=6.05 $Y=0.675 $X2=0
+ $Y2=0
cc_979 N_A_659_113#_c_911_n N_VGND_c_2836_n 0.0150383f $X=6.135 $Y=0.34 $X2=0
+ $Y2=0
cc_980 N_A_659_113#_c_910_n N_VGND_c_2837_n 0.0122839f $X=6.725 $Y=0.34 $X2=0
+ $Y2=0
cc_981 N_A_659_113#_c_912_n N_VGND_c_2837_n 0.00727799f $X=6.81 $Y=1.13 $X2=0
+ $Y2=0
cc_982 N_A_659_113#_c_913_n N_VGND_c_2837_n 0.0202823f $X=7.535 $Y=1.215 $X2=0
+ $Y2=0
cc_983 N_A_659_113#_c_915_n N_VGND_c_2837_n 0.0281254f $X=7.62 $Y=1.13 $X2=0
+ $Y2=0
cc_984 N_A_659_113#_c_917_n N_VGND_c_2837_n 0.0147457f $X=7.705 $Y=0.34 $X2=0
+ $Y2=0
cc_985 N_A_659_113#_c_916_n N_VGND_c_2838_n 0.00607851f $X=10.085 $Y=0.34 $X2=0
+ $Y2=0
cc_986 N_A_659_113#_c_918_n N_VGND_c_2838_n 0.0052832f $X=10.17 $Y=1.545 $X2=0
+ $Y2=0
cc_987 N_A_659_113#_c_907_n N_VGND_c_2845_n 0.00283604f $X=5.965 $Y=0.76 $X2=0
+ $Y2=0
cc_988 N_A_659_113#_c_910_n N_VGND_c_2845_n 0.0501353f $X=6.725 $Y=0.34 $X2=0
+ $Y2=0
cc_989 N_A_659_113#_c_911_n N_VGND_c_2845_n 0.0120568f $X=6.135 $Y=0.34 $X2=0
+ $Y2=0
cc_990 N_A_659_113#_c_896_n N_VGND_c_2850_n 0.00324627f $X=3.37 $Y=1.225 $X2=0
+ $Y2=0
cc_991 N_A_659_113#_c_908_n N_VGND_c_2850_n 2.37437e-19 $X=5.78 $Y=0.76 $X2=0
+ $Y2=0
cc_992 N_A_659_113#_c_916_n N_VGND_c_2851_n 0.164795f $X=10.085 $Y=0.34 $X2=0
+ $Y2=0
cc_993 N_A_659_113#_c_917_n N_VGND_c_2851_n 0.0115893f $X=7.705 $Y=0.34 $X2=0
+ $Y2=0
cc_994 N_A_659_113#_c_896_n N_VGND_c_2854_n 0.00375425f $X=3.37 $Y=1.225 $X2=0
+ $Y2=0
cc_995 N_A_659_113#_c_907_n N_VGND_c_2854_n 0.00480001f $X=5.965 $Y=0.76 $X2=0
+ $Y2=0
cc_996 N_A_659_113#_c_908_n N_VGND_c_2854_n 0.00188442f $X=5.78 $Y=0.76 $X2=0
+ $Y2=0
cc_997 N_A_659_113#_c_910_n N_VGND_c_2854_n 0.0287839f $X=6.725 $Y=0.34 $X2=0
+ $Y2=0
cc_998 N_A_659_113#_c_911_n N_VGND_c_2854_n 0.00658475f $X=6.135 $Y=0.34 $X2=0
+ $Y2=0
cc_999 N_A_659_113#_c_916_n N_VGND_c_2854_n 0.0858223f $X=10.085 $Y=0.34 $X2=0
+ $Y2=0
cc_1000 N_A_659_113#_c_917_n N_VGND_c_2854_n 0.00583135f $X=7.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1001 N_A_659_113#_c_912_n A_1336_97# 0.00223521f $X=6.81 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_1002 N_A_659_113#_c_918_n A_2002_125# 0.00557298f $X=10.17 $Y=1.545 $X2=-0.19
+ $Y2=-0.245
cc_1003 N_A_659_113#_c_918_n N_A_2074_125#_c_3022_n 0.0269936f $X=10.17 $Y=1.545
+ $X2=0 $Y2=0
cc_1004 N_A_659_113#_c_919_n N_A_2074_125#_c_3023_n 0.0661397f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_1005 N_A_659_113#_c_918_n N_A_2074_125#_c_3024_n 0.0137141f $X=10.17 $Y=1.545
+ $X2=0 $Y2=0
cc_1006 N_A_659_113#_c_919_n N_A_2074_125#_c_3024_n 0.0137141f $X=12.505 $Y=1.63
+ $X2=0 $Y2=0
cc_1007 N_A_659_113#_c_923_n A_3056_72# 0.00130185f $X=15.405 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_1008 N_A_1068_21#_M1035_g N_A_887_139#_M1009_g 0.0160317f $X=5.975 $Y=2.885
+ $X2=0 $Y2=0
cc_1009 N_A_1068_21#_c_1256_n N_A_887_139#_M1009_g 0.0113581f $X=6.68 $Y=2.375
+ $X2=0 $Y2=0
cc_1010 N_A_1068_21#_c_1257_n N_A_887_139#_M1009_g 0.0242435f $X=6.065 $Y=2.35
+ $X2=0 $Y2=0
cc_1011 N_A_1068_21#_c_1259_n N_A_887_139#_M1009_g 0.0054957f $X=6.845 $Y=2.375
+ $X2=0 $Y2=0
cc_1012 N_A_1068_21#_c_1251_n N_A_887_139#_M1038_g 0.0263737f $X=6.155 $Y=1.345
+ $X2=0 $Y2=0
cc_1013 N_A_1068_21#_c_1252_n N_A_887_139#_M1038_g 0.00577587f $X=6.305 $Y=1.157
+ $X2=0 $Y2=0
cc_1014 N_A_1068_21#_c_1253_n N_A_887_139#_M1038_g 0.00577329f $X=6.39 $Y=0.76
+ $X2=0 $Y2=0
cc_1015 N_A_1068_21#_c_1254_n N_A_887_139#_M1038_g 0.0185068f $X=6.065 $Y=2.185
+ $X2=0 $Y2=0
cc_1016 N_A_1068_21#_c_1257_n N_A_887_139#_c_1354_n 0.00274379f $X=6.065 $Y=2.35
+ $X2=0 $Y2=0
cc_1017 N_A_1068_21#_c_1258_n N_A_887_139#_c_1354_n 0.0102135f $X=6.23 $Y=2.365
+ $X2=0 $Y2=0
cc_1018 N_A_1068_21#_c_1254_n N_A_887_139#_c_1354_n 4.97396e-19 $X=6.065
+ $Y=2.185 $X2=0 $Y2=0
cc_1019 N_A_1068_21#_c_1256_n N_A_887_139#_c_1355_n 0.0171186f $X=6.68 $Y=2.375
+ $X2=0 $Y2=0
cc_1020 N_A_1068_21#_c_1254_n N_A_887_139#_c_1355_n 7.45832e-19 $X=6.065
+ $Y=2.185 $X2=0 $Y2=0
cc_1021 N_A_1068_21#_c_1256_n N_A_887_139#_c_1356_n 0.00238453f $X=6.68 $Y=2.375
+ $X2=0 $Y2=0
cc_1022 N_A_1068_21#_c_1259_n N_A_887_139#_c_1356_n 0.00204323f $X=6.845
+ $Y=2.375 $X2=0 $Y2=0
cc_1023 N_A_1068_21#_c_1254_n N_A_887_139#_c_1356_n 0.0242435f $X=6.065 $Y=2.185
+ $X2=0 $Y2=0
cc_1024 N_A_1068_21#_c_1259_n N_A_887_139#_c_1357_n 0.0236172f $X=6.845 $Y=2.375
+ $X2=0 $Y2=0
cc_1025 N_A_1068_21#_c_1256_n N_A_887_139#_c_1360_n 0.014358f $X=6.68 $Y=2.375
+ $X2=0 $Y2=0
cc_1026 N_A_1068_21#_c_1257_n N_A_887_139#_c_1360_n 0.00496257f $X=6.065 $Y=2.35
+ $X2=0 $Y2=0
cc_1027 N_A_1068_21#_c_1258_n N_A_887_139#_c_1360_n 0.0230706f $X=6.23 $Y=2.365
+ $X2=0 $Y2=0
cc_1028 N_A_1068_21#_c_1254_n N_A_887_139#_c_1360_n 0.0110711f $X=6.065 $Y=2.185
+ $X2=0 $Y2=0
cc_1029 N_A_1068_21#_c_1259_n N_SET_B_M1027_g 0.00616886f $X=6.845 $Y=2.375
+ $X2=0 $Y2=0
cc_1030 N_A_1068_21#_M1035_g N_VPWR_c_2357_n 0.0121054f $X=5.975 $Y=2.885 $X2=0
+ $Y2=0
cc_1031 N_A_1068_21#_c_1257_n N_VPWR_c_2357_n 0.00495888f $X=6.065 $Y=2.35 $X2=0
+ $Y2=0
cc_1032 N_A_1068_21#_c_1258_n N_VPWR_c_2357_n 0.0251627f $X=6.23 $Y=2.365 $X2=0
+ $Y2=0
cc_1033 N_A_1068_21#_c_1259_n N_VPWR_c_2357_n 0.00176295f $X=6.845 $Y=2.375
+ $X2=0 $Y2=0
cc_1034 N_A_1068_21#_c_1259_n N_VPWR_c_2358_n 0.025384f $X=6.845 $Y=2.375 $X2=0
+ $Y2=0
cc_1035 N_A_1068_21#_M1035_g N_VPWR_c_2360_n 0.00486043f $X=5.975 $Y=2.885 $X2=0
+ $Y2=0
cc_1036 N_A_1068_21#_c_1259_n N_VPWR_c_2364_n 0.00609883f $X=6.845 $Y=2.375
+ $X2=0 $Y2=0
cc_1037 N_A_1068_21#_M1009_d N_VPWR_c_2354_n 0.00181679f $X=6.59 $Y=2.675 $X2=0
+ $Y2=0
cc_1038 N_A_1068_21#_M1035_g N_VPWR_c_2354_n 0.00337932f $X=5.975 $Y=2.885 $X2=0
+ $Y2=0
cc_1039 N_A_1068_21#_c_1259_n N_VPWR_c_2354_n 9.62626e-19 $X=6.845 $Y=2.375
+ $X2=0 $Y2=0
cc_1040 N_A_1068_21#_M1009_d N_KAPWR_c_2677_n 0.00251772f $X=6.59 $Y=2.675 $X2=0
+ $Y2=0
cc_1041 N_A_1068_21#_M1035_g N_KAPWR_c_2677_n 0.00365667f $X=5.975 $Y=2.885
+ $X2=0 $Y2=0
cc_1042 N_A_1068_21#_c_1256_n N_KAPWR_c_2677_n 0.0147164f $X=6.68 $Y=2.375 $X2=0
+ $Y2=0
cc_1043 N_A_1068_21#_c_1258_n N_KAPWR_c_2677_n 0.0075243f $X=6.23 $Y=2.365 $X2=0
+ $Y2=0
cc_1044 N_A_1068_21#_c_1259_n N_KAPWR_c_2677_n 0.01347f $X=6.845 $Y=2.375 $X2=0
+ $Y2=0
cc_1045 N_A_1068_21#_c_1248_n N_VGND_c_2836_n 0.00919702f $X=5.415 $Y=0.765
+ $X2=0 $Y2=0
cc_1046 N_A_1068_21#_c_1249_n N_VGND_c_2836_n 0.00177054f $X=5.99 $Y=0.84 $X2=0
+ $Y2=0
cc_1047 N_A_1068_21#_c_1249_n N_VGND_c_2845_n 9.19576e-19 $X=5.99 $Y=0.84 $X2=0
+ $Y2=0
cc_1048 N_A_1068_21#_c_1248_n N_VGND_c_2850_n 0.00471611f $X=5.415 $Y=0.765
+ $X2=0 $Y2=0
cc_1049 N_A_1068_21#_c_1248_n N_VGND_c_2854_n 0.00805858f $X=5.415 $Y=0.765
+ $X2=0 $Y2=0
cc_1050 N_A_887_139#_M1038_g N_SET_B_M1003_g 0.0520937f $X=6.605 $Y=0.695 $X2=0
+ $Y2=0
cc_1051 N_A_887_139#_M1040_g N_SET_B_M1003_g 0.0165171f $X=7.63 $Y=0.945 $X2=0
+ $Y2=0
cc_1052 N_A_887_139#_M1009_g N_SET_B_M1027_g 0.0160548f $X=6.515 $Y=2.885 $X2=0
+ $Y2=0
cc_1053 N_A_887_139#_M1038_g N_SET_B_M1027_g 0.0118921f $X=6.605 $Y=0.695 $X2=0
+ $Y2=0
cc_1054 N_A_887_139#_M1032_g N_SET_B_M1027_g 0.013597f $X=7.63 $Y=2.675 $X2=0
+ $Y2=0
cc_1055 N_A_887_139#_c_1356_n N_SET_B_M1027_g 0.0209878f $X=6.605 $Y=1.93 $X2=0
+ $Y2=0
cc_1056 N_A_887_139#_c_1357_n N_SET_B_M1027_g 0.0147384f $X=7.51 $Y=1.93 $X2=0
+ $Y2=0
cc_1057 N_A_887_139#_c_1346_n N_SET_B_M1027_g 0.0327128f $X=7.51 $Y=1.93 $X2=0
+ $Y2=0
cc_1058 N_A_887_139#_M1040_g N_SET_B_c_2001_n 0.00825762f $X=7.63 $Y=0.945 $X2=0
+ $Y2=0
cc_1059 N_A_887_139#_M1040_g N_SET_B_c_2008_n 0.00814335f $X=7.63 $Y=0.945 $X2=0
+ $Y2=0
cc_1060 N_A_887_139#_c_1357_n N_SET_B_c_2008_n 3.01859e-19 $X=7.51 $Y=1.93 $X2=0
+ $Y2=0
cc_1061 N_A_887_139#_M1009_g N_VPWR_c_2357_n 0.0126704f $X=6.515 $Y=2.885 $X2=0
+ $Y2=0
cc_1062 N_A_887_139#_c_1354_n N_VPWR_c_2357_n 0.00910813f $X=5.37 $Y=2.865 $X2=0
+ $Y2=0
cc_1063 N_A_887_139#_M1009_g N_VPWR_c_2358_n 0.00658944f $X=6.515 $Y=2.885 $X2=0
+ $Y2=0
cc_1064 N_A_887_139#_M1032_g N_VPWR_c_2358_n 0.0177078f $X=7.63 $Y=2.675 $X2=0
+ $Y2=0
cc_1065 N_A_887_139#_c_1357_n N_VPWR_c_2358_n 0.023879f $X=7.51 $Y=1.93 $X2=0
+ $Y2=0
cc_1066 N_A_887_139#_c_1346_n N_VPWR_c_2358_n 0.00511968f $X=7.51 $Y=1.93 $X2=0
+ $Y2=0
cc_1067 N_A_887_139#_c_1354_n N_VPWR_c_2360_n 0.018989f $X=5.37 $Y=2.865 $X2=0
+ $Y2=0
cc_1068 N_A_887_139#_M1009_g N_VPWR_c_2364_n 0.00585385f $X=6.515 $Y=2.885 $X2=0
+ $Y2=0
cc_1069 N_A_887_139#_M1032_g N_VPWR_c_2365_n 0.00486043f $X=7.63 $Y=2.675 $X2=0
+ $Y2=0
cc_1070 N_A_887_139#_M1005_d N_VPWR_c_2354_n 0.00114239f $X=5.23 $Y=2.675 $X2=0
+ $Y2=0
cc_1071 N_A_887_139#_M1009_g N_VPWR_c_2354_n 0.00680348f $X=6.515 $Y=2.885 $X2=0
+ $Y2=0
cc_1072 N_A_887_139#_M1032_g N_VPWR_c_2354_n 0.00446301f $X=7.63 $Y=2.675 $X2=0
+ $Y2=0
cc_1073 N_A_887_139#_c_1354_n N_VPWR_c_2354_n 0.00303042f $X=5.37 $Y=2.865 $X2=0
+ $Y2=0
cc_1074 N_A_887_139#_c_1345_n N_A_189_119#_c_2520_n 0.00749985f $X=4.855
+ $Y=1.905 $X2=0 $Y2=0
cc_1075 N_A_887_139#_c_1347_n N_A_189_119#_c_2520_n 0.0153706f $X=4.855 $Y=0.905
+ $X2=0 $Y2=0
cc_1076 N_A_887_139#_c_1345_n N_A_189_119#_c_2521_n 0.0142489f $X=4.855 $Y=1.905
+ $X2=0 $Y2=0
cc_1077 N_A_887_139#_c_1347_n N_A_189_119#_c_2521_n 0.0128425f $X=4.855 $Y=0.905
+ $X2=0 $Y2=0
cc_1078 N_A_887_139#_c_1345_n N_A_189_119#_c_2523_n 0.0262798f $X=4.855 $Y=1.905
+ $X2=0 $Y2=0
cc_1079 N_A_887_139#_c_1352_n N_A_189_119#_c_2523_n 0.00262249f $X=5.205 $Y=1.99
+ $X2=0 $Y2=0
cc_1080 N_A_887_139#_c_1353_n N_A_189_119#_c_2523_n 0.0194251f $X=4.94 $Y=1.99
+ $X2=0 $Y2=0
cc_1081 N_A_887_139#_c_1354_n N_A_189_119#_c_2523_n 0.0371074f $X=5.37 $Y=2.865
+ $X2=0 $Y2=0
cc_1082 N_A_887_139#_M1040_g N_A_1541_125#_c_2636_n 0.00362071f $X=7.63 $Y=0.945
+ $X2=0 $Y2=0
cc_1083 N_A_887_139#_M1040_g N_A_1541_125#_c_2637_n 0.00104849f $X=7.63 $Y=0.945
+ $X2=0 $Y2=0
cc_1084 N_A_887_139#_M1040_g N_A_1541_125#_c_2653_n 8.1802e-19 $X=7.63 $Y=0.945
+ $X2=0 $Y2=0
cc_1085 N_A_887_139#_M1009_g N_KAPWR_c_2677_n 0.00948585f $X=6.515 $Y=2.885
+ $X2=0 $Y2=0
cc_1086 N_A_887_139#_M1032_g N_KAPWR_c_2677_n 0.00688162f $X=7.63 $Y=2.675 $X2=0
+ $Y2=0
cc_1087 N_A_887_139#_c_1352_n N_KAPWR_c_2677_n 0.00559514f $X=5.205 $Y=1.99
+ $X2=0 $Y2=0
cc_1088 N_A_887_139#_c_1353_n N_KAPWR_c_2677_n 0.00125303f $X=4.94 $Y=1.99 $X2=0
+ $Y2=0
cc_1089 N_A_887_139#_c_1354_n N_KAPWR_c_2677_n 0.0390621f $X=5.37 $Y=2.865 $X2=0
+ $Y2=0
cc_1090 N_A_887_139#_c_1355_n N_KAPWR_c_2677_n 3.34088e-19 $X=6.582 $Y=1.952
+ $X2=0 $Y2=0
cc_1091 N_A_887_139#_c_1357_n N_KAPWR_c_2677_n 0.0122846f $X=7.51 $Y=1.93 $X2=0
+ $Y2=0
cc_1092 N_A_887_139#_c_1360_n N_KAPWR_c_2677_n 0.0110982f $X=6.44 $Y=1.952 $X2=0
+ $Y2=0
cc_1093 N_A_887_139#_M1040_g N_VGND_c_2837_n 0.00174045f $X=7.63 $Y=0.945 $X2=0
+ $Y2=0
cc_1094 N_A_887_139#_M1038_g N_VGND_c_2845_n 7.35405e-19 $X=6.605 $Y=0.695 $X2=0
+ $Y2=0
cc_1095 N_A_1972_99#_M1006_g N_A_2216_99#_c_1617_n 0.00119631f $X=10.295
+ $Y=0.835 $X2=0 $Y2=0
cc_1096 N_A_1972_99#_c_1531_n N_A_2216_99#_c_1618_n 4.8095e-19 $X=12.93 $Y=1.1
+ $X2=0 $Y2=0
cc_1097 N_A_1972_99#_c_1481_n N_A_2216_99#_c_1618_n 0.0148351f $X=14.425
+ $Y=1.325 $X2=0 $Y2=0
cc_1098 N_A_1972_99#_c_1489_n N_A_2216_99#_M1024_g 0.00497567f $X=12.845 $Y=1.97
+ $X2=0 $Y2=0
cc_1099 N_A_1972_99#_c_1480_n N_A_2216_99#_M1024_g 0.00923332f $X=12.93 $Y=1.885
+ $X2=0 $Y2=0
cc_1100 N_A_1972_99#_c_1481_n N_A_2216_99#_M1024_g 0.0111549f $X=14.425 $Y=1.325
+ $X2=0 $Y2=0
cc_1101 N_A_1972_99#_c_1531_n N_A_2216_99#_c_1620_n 0.00343408f $X=12.93 $Y=1.1
+ $X2=0 $Y2=0
cc_1102 N_A_1972_99#_c_1488_n N_A_1728_125#_c_1791_n 0.00945214f $X=11.475
+ $Y=1.97 $X2=0 $Y2=0
cc_1103 N_A_1972_99#_c_1491_n N_A_1728_125#_c_1791_n 6.01453e-19 $X=10.82
+ $Y=1.97 $X2=0 $Y2=0
cc_1104 N_A_1972_99#_c_1493_n N_A_1728_125#_c_1791_n 0.00598118f $X=11.64
+ $Y=1.97 $X2=0 $Y2=0
cc_1105 N_A_1972_99#_c_1488_n N_A_1728_125#_c_1792_n 0.00113446f $X=11.475
+ $Y=1.97 $X2=0 $Y2=0
cc_1106 N_A_1972_99#_c_1489_n N_A_1728_125#_c_1792_n 0.00970206f $X=12.845
+ $Y=1.97 $X2=0 $Y2=0
cc_1107 N_A_1972_99#_c_1493_n N_A_1728_125#_c_1792_n 0.00990994f $X=11.64
+ $Y=1.97 $X2=0 $Y2=0
cc_1108 N_A_1972_99#_c_1488_n N_A_1728_125#_c_1793_n 0.00150381f $X=11.475
+ $Y=1.97 $X2=0 $Y2=0
cc_1109 N_A_1972_99#_c_1492_n N_A_1728_125#_c_1793_n 0.0175613f $X=10.82 $Y=2.05
+ $X2=0 $Y2=0
cc_1110 N_A_1972_99#_c_1485_n N_A_1728_125#_c_1793_n 0.00556646f $X=10.82
+ $Y=1.885 $X2=0 $Y2=0
cc_1111 N_A_1972_99#_c_1489_n N_A_1728_125#_c_1795_n 0.0131414f $X=12.845
+ $Y=1.97 $X2=0 $Y2=0
cc_1112 N_A_1972_99#_c_1493_n N_A_1728_125#_c_1795_n 0.00488109f $X=11.64
+ $Y=1.97 $X2=0 $Y2=0
cc_1113 N_A_1972_99#_c_1531_n N_A_1728_125#_M1041_g 0.00268644f $X=12.93 $Y=1.1
+ $X2=0 $Y2=0
cc_1114 N_A_1972_99#_c_1480_n N_A_1728_125#_M1041_g 0.00534166f $X=12.93
+ $Y=1.885 $X2=0 $Y2=0
cc_1115 N_A_1972_99#_c_1482_n N_A_1728_125#_M1041_g 0.00131304f $X=12.93
+ $Y=1.325 $X2=0 $Y2=0
cc_1116 N_A_1972_99#_c_1489_n N_A_1728_125#_c_1799_n 0.0103612f $X=12.845
+ $Y=1.97 $X2=0 $Y2=0
cc_1117 N_A_1972_99#_M1018_s N_A_1728_125#_c_1801_n 0.0132055f $X=11.495
+ $Y=2.005 $X2=0 $Y2=0
cc_1118 N_A_1972_99#_c_1486_n N_A_1728_125#_c_1802_n 0.0215439f $X=14.705
+ $Y=2.065 $X2=0 $Y2=0
cc_1119 N_A_1972_99#_c_1486_n N_A_1728_125#_c_1844_n 0.00122227f $X=14.705
+ $Y=2.065 $X2=0 $Y2=0
cc_1120 N_A_1972_99#_c_1486_n N_A_1728_125#_c_1849_n 0.00467643f $X=14.705
+ $Y=2.065 $X2=0 $Y2=0
cc_1121 N_A_1972_99#_M1046_g N_SET_B_c_2001_n 0.00737859f $X=9.935 $Y=0.835
+ $X2=0 $Y2=0
cc_1122 N_A_1972_99#_M1006_g N_SET_B_c_2001_n 0.00888494f $X=10.295 $Y=0.835
+ $X2=0 $Y2=0
cc_1123 N_A_1972_99#_M1006_g N_SET_B_M1008_g 0.0107281f $X=10.295 $Y=0.835 $X2=0
+ $Y2=0
cc_1124 N_A_1972_99#_c_1477_n N_SET_B_M1008_g 0.00773791f $X=10.655 $Y=1.5 $X2=0
+ $Y2=0
cc_1125 N_A_1972_99#_c_1481_n N_SET_B_c_2005_n 0.0119548f $X=14.425 $Y=1.325
+ $X2=0 $Y2=0
cc_1126 N_A_1972_99#_c_1481_n N_SET_B_c_2006_n 0.00320674f $X=14.425 $Y=1.325
+ $X2=0 $Y2=0
cc_1127 N_A_1972_99#_c_1483_n N_SET_B_c_2007_n 0.00130453f $X=14.59 $Y=1.205
+ $X2=0 $Y2=0
cc_1128 N_A_1972_99#_c_1484_n N_SET_B_c_2007_n 0.020195f $X=14.59 $Y=1.205 $X2=0
+ $Y2=0
cc_1129 N_A_1972_99#_c_1480_n SET_B 0.00884665f $X=12.93 $Y=1.885 $X2=0 $Y2=0
cc_1130 N_A_1972_99#_c_1481_n SET_B 0.0237746f $X=14.425 $Y=1.325 $X2=0 $Y2=0
cc_1131 N_A_1972_99#_c_1481_n N_SET_B_c_2011_n 0.00124763f $X=14.425 $Y=1.325
+ $X2=0 $Y2=0
cc_1132 N_A_1972_99#_c_1481_n N_SET_B_c_2012_n 0.00530439f $X=14.425 $Y=1.325
+ $X2=0 $Y2=0
cc_1133 N_A_1972_99#_c_1484_n N_SET_B_c_2012_n 4.08455e-19 $X=14.59 $Y=1.205
+ $X2=0 $Y2=0
cc_1134 N_A_1972_99#_c_1483_n N_CLK_M1015_g 7.21666e-19 $X=14.59 $Y=1.205 $X2=0
+ $Y2=0
cc_1135 N_A_1972_99#_c_1484_n N_CLK_M1015_g 0.00902742f $X=14.59 $Y=1.205 $X2=0
+ $Y2=0
cc_1136 N_A_1972_99#_c_1486_n N_CLK_M1039_g 0.0185829f $X=14.705 $Y=2.065 $X2=0
+ $Y2=0
cc_1137 N_A_1972_99#_c_1479_n N_CLK_M1039_g 0.00335298f $X=14.705 $Y=1.94 $X2=0
+ $Y2=0
cc_1138 N_A_1972_99#_c_1486_n CLK 0.00554066f $X=14.705 $Y=2.065 $X2=0 $Y2=0
cc_1139 N_A_1972_99#_c_1479_n CLK 0.00364869f $X=14.705 $Y=1.94 $X2=0 $Y2=0
cc_1140 N_A_1972_99#_c_1483_n CLK 0.0149975f $X=14.59 $Y=1.205 $X2=0 $Y2=0
cc_1141 N_A_1972_99#_c_1484_n CLK 0.00298489f $X=14.59 $Y=1.205 $X2=0 $Y2=0
cc_1142 N_A_1972_99#_c_1483_n N_CLK_c_2123_n 2.43687e-19 $X=14.59 $Y=1.205 $X2=0
+ $Y2=0
cc_1143 N_A_1972_99#_c_1484_n N_CLK_c_2123_n 0.0214809f $X=14.59 $Y=1.205 $X2=0
+ $Y2=0
cc_1144 N_A_1972_99#_c_1486_n N_VPWR_c_2365_n 0.00569155f $X=14.705 $Y=2.065
+ $X2=0 $Y2=0
cc_1145 N_A_1972_99#_c_1486_n N_VPWR_c_2354_n 0.00781321f $X=14.705 $Y=2.065
+ $X2=0 $Y2=0
cc_1146 N_A_1972_99#_c_1489_n N_KAPWR_M1018_d 0.0020475f $X=12.845 $Y=1.97
+ $X2=-0.19 $Y2=-0.245
cc_1147 N_A_1972_99#_c_1486_n N_KAPWR_c_2675_n 0.0143859f $X=14.705 $Y=2.065
+ $X2=0 $Y2=0
cc_1148 N_A_1972_99#_M1018_s N_KAPWR_c_2677_n 0.00672939f $X=11.495 $Y=2.005
+ $X2=0 $Y2=0
cc_1149 N_A_1972_99#_c_1486_n N_KAPWR_c_2677_n 0.0087779f $X=14.705 $Y=2.065
+ $X2=0 $Y2=0
cc_1150 N_A_1972_99#_c_1486_n N_KAPWR_c_2678_n 0.00951242f $X=14.705 $Y=2.065
+ $X2=0 $Y2=0
cc_1151 N_A_1972_99#_M1006_g N_VGND_c_2838_n 4.52274e-19 $X=10.295 $Y=0.835
+ $X2=0 $Y2=0
cc_1152 N_A_1972_99#_M1006_g N_VGND_c_2854_n 7.30987e-19 $X=10.295 $Y=0.835
+ $X2=0 $Y2=0
cc_1153 N_A_1972_99#_M1006_g N_A_2074_125#_c_3022_n 0.00151769f $X=10.295
+ $Y=0.835 $X2=0 $Y2=0
cc_1154 N_A_1972_99#_c_1477_n N_A_2074_125#_c_3023_n 0.00259696f $X=10.655
+ $Y=1.5 $X2=0 $Y2=0
cc_1155 N_A_1972_99#_M1006_g N_A_2074_125#_c_3024_n 0.00289461f $X=10.295
+ $Y=0.835 $X2=0 $Y2=0
cc_1156 N_A_1972_99#_c_1477_n N_A_2074_125#_c_3024_n 0.00394113f $X=10.655
+ $Y=1.5 $X2=0 $Y2=0
cc_1157 N_A_2216_99#_c_1622_n N_A_1728_125#_c_1792_n 0.0116887f $X=11.79 $Y=1.29
+ $X2=0 $Y2=0
cc_1158 N_A_2216_99#_c_1634_n N_A_1728_125#_c_1792_n 0.00421114f $X=11.625
+ $Y=1.29 $X2=0 $Y2=0
cc_1159 N_A_2216_99#_c_1617_n N_A_1728_125#_c_1793_n 0.00421114f $X=11.23
+ $Y=1.23 $X2=0 $Y2=0
cc_1160 N_A_2216_99#_c_1621_n N_A_1728_125#_M1051_g 0.00837911f $X=12.165
+ $Y=1.25 $X2=0 $Y2=0
cc_1161 N_A_2216_99#_c_1622_n N_A_1728_125#_M1051_g 0.021569f $X=11.79 $Y=1.29
+ $X2=0 $Y2=0
cc_1162 N_A_2216_99#_c_1623_n N_A_1728_125#_M1051_g 0.0202641f $X=12.25 $Y=1.125
+ $X2=0 $Y2=0
cc_1163 N_A_2216_99#_M1024_g N_A_1728_125#_c_1795_n 0.0340147f $X=13.165 $Y=2.57
+ $X2=0 $Y2=0
cc_1164 N_A_2216_99#_c_1618_n N_A_1728_125#_M1041_g 0.00977699f $X=13.165
+ $Y=1.37 $X2=0 $Y2=0
cc_1165 N_A_2216_99#_c_1621_n N_A_1728_125#_M1041_g 9.04319e-19 $X=12.165
+ $Y=1.25 $X2=0 $Y2=0
cc_1166 N_A_2216_99#_c_1623_n N_A_1728_125#_M1041_g 0.00310851f $X=12.25
+ $Y=1.125 $X2=0 $Y2=0
cc_1167 N_A_2216_99#_c_1624_n N_A_1728_125#_M1041_g 0.00114816f $X=13.525
+ $Y=0.34 $X2=0 $Y2=0
cc_1168 N_A_2216_99#_c_1633_n N_A_1728_125#_M1041_g 0.0104189f $X=13.69 $Y=0.63
+ $X2=0 $Y2=0
cc_1169 N_A_2216_99#_c_1631_n N_A_1728_125#_c_1784_n 0.00456942f $X=16.67
+ $Y=2.065 $X2=0 $Y2=0
cc_1170 N_A_2216_99#_c_1630_n N_A_1728_125#_c_1786_n 0.00274791f $X=16.645
+ $Y=1.05 $X2=0 $Y2=0
cc_1171 N_A_2216_99#_c_1630_n N_A_1728_125#_M1007_g 0.00115212f $X=16.645
+ $Y=1.05 $X2=0 $Y2=0
cc_1172 N_A_2216_99#_M1024_g N_A_1728_125#_c_1799_n 0.00786837f $X=13.165
+ $Y=2.57 $X2=0 $Y2=0
cc_1173 N_A_2216_99#_M1024_g N_A_1728_125#_c_1830_n 0.0137296f $X=13.165 $Y=2.57
+ $X2=0 $Y2=0
cc_1174 N_A_2216_99#_M1045_d N_A_1728_125#_c_1802_n 0.0063993f $X=16.53 $Y=1.92
+ $X2=0 $Y2=0
cc_1175 N_A_2216_99#_c_1631_n N_A_1728_125#_c_1802_n 0.0248434f $X=16.67
+ $Y=2.065 $X2=0 $Y2=0
cc_1176 N_A_2216_99#_c_1631_n N_A_1728_125#_c_1803_n 0.0220759f $X=16.67
+ $Y=2.065 $X2=0 $Y2=0
cc_1177 N_A_2216_99#_M1024_g N_A_1728_125#_c_1805_n 0.00125309f $X=13.165
+ $Y=2.57 $X2=0 $Y2=0
cc_1178 N_A_2216_99#_c_1631_n N_A_1728_125#_c_1789_n 0.0264121f $X=16.67
+ $Y=2.065 $X2=0 $Y2=0
cc_1179 N_A_2216_99#_c_1630_n N_A_1728_125#_c_1790_n 0.00164886f $X=16.645
+ $Y=1.05 $X2=0 $Y2=0
cc_1180 N_A_2216_99#_c_1631_n N_A_1728_125#_c_1790_n 0.00342519f $X=16.67
+ $Y=2.065 $X2=0 $Y2=0
cc_1181 N_A_2216_99#_c_1616_n N_SET_B_M1008_g 0.0118531f $X=11.155 $Y=1.155
+ $X2=0 $Y2=0
cc_1182 N_A_2216_99#_c_1616_n N_SET_B_c_2004_n 0.00895007f $X=11.155 $Y=1.155
+ $X2=0 $Y2=0
cc_1183 N_A_2216_99#_c_1624_n N_SET_B_c_2004_n 0.0220144f $X=13.525 $Y=0.34
+ $X2=0 $Y2=0
cc_1184 N_A_2216_99#_c_1625_n N_SET_B_c_2004_n 0.00169616f $X=12.335 $Y=0.34
+ $X2=0 $Y2=0
cc_1185 N_A_2216_99#_c_1626_n N_SET_B_c_2004_n 0.00281801f $X=15.745 $Y=0.34
+ $X2=0 $Y2=0
cc_1186 N_A_2216_99#_c_1632_n N_SET_B_c_2004_n 0.00249866f $X=13.69 $Y=0.34
+ $X2=0 $Y2=0
cc_1187 N_A_2216_99#_c_1633_n N_SET_B_c_2004_n 0.033182f $X=13.69 $Y=0.63 $X2=0
+ $Y2=0
cc_1188 N_A_2216_99#_M1024_g N_SET_B_M1043_g 0.0723548f $X=13.165 $Y=2.57 $X2=0
+ $Y2=0
cc_1189 N_A_2216_99#_c_1620_n N_SET_B_c_2006_n 0.00600446f $X=13.395 $Y=1.22
+ $X2=0 $Y2=0
cc_1190 N_A_2216_99#_c_1633_n N_SET_B_c_2006_n 0.00437137f $X=13.69 $Y=0.63
+ $X2=0 $Y2=0
cc_1191 N_A_2216_99#_c_1620_n N_SET_B_c_2007_n 0.0052695f $X=13.395 $Y=1.22
+ $X2=0 $Y2=0
cc_1192 N_A_2216_99#_c_1626_n N_SET_B_c_2007_n 0.0115145f $X=15.745 $Y=0.34
+ $X2=0 $Y2=0
cc_1193 N_A_2216_99#_c_1632_n N_SET_B_c_2007_n 0.00308445f $X=13.69 $Y=0.34
+ $X2=0 $Y2=0
cc_1194 N_A_2216_99#_c_1633_n N_SET_B_c_2007_n 0.0211089f $X=13.69 $Y=0.63 $X2=0
+ $Y2=0
cc_1195 N_A_2216_99#_M1024_g SET_B 0.00103858f $X=13.165 $Y=2.57 $X2=0 $Y2=0
cc_1196 N_A_2216_99#_M1024_g N_SET_B_c_2011_n 0.0218424f $X=13.165 $Y=2.57 $X2=0
+ $Y2=0
cc_1197 N_A_2216_99#_c_1618_n N_SET_B_c_2012_n 0.00600446f $X=13.165 $Y=1.37
+ $X2=0 $Y2=0
cc_1198 N_A_2216_99#_M1024_g N_SET_B_c_2012_n 0.00709514f $X=13.165 $Y=2.57
+ $X2=0 $Y2=0
cc_1199 N_A_2216_99#_c_1626_n N_CLK_M1015_g 0.010978f $X=15.745 $Y=0.34 $X2=0
+ $Y2=0
cc_1200 N_A_2216_99#_c_1626_n N_SLEEP_B_M1014_g 0.011362f $X=15.745 $Y=0.34
+ $X2=0 $Y2=0
cc_1201 N_A_2216_99#_c_1627_n N_SLEEP_B_M1014_g 0.0054219f $X=15.83 $Y=0.88
+ $X2=0 $Y2=0
cc_1202 N_A_2216_99#_c_1629_n N_SLEEP_B_M1014_g 5.08826e-19 $X=15.915 $Y=0.965
+ $X2=0 $Y2=0
cc_1203 N_A_2216_99#_c_1626_n N_SLEEP_B_M1049_g 0.00359132f $X=15.745 $Y=0.34
+ $X2=0 $Y2=0
cc_1204 N_A_2216_99#_c_1627_n N_SLEEP_B_M1049_g 0.00850129f $X=15.83 $Y=0.88
+ $X2=0 $Y2=0
cc_1205 N_A_2216_99#_c_1628_n N_SLEEP_B_M1049_g 0.00653163f $X=16.455 $Y=0.965
+ $X2=0 $Y2=0
cc_1206 N_A_2216_99#_c_1629_n N_SLEEP_B_M1049_g 6.34888e-19 $X=15.915 $Y=0.965
+ $X2=0 $Y2=0
cc_1207 N_A_2216_99#_c_1631_n N_SLEEP_B_c_2171_n 0.00911871f $X=16.67 $Y=2.065
+ $X2=0 $Y2=0
cc_1208 N_A_2216_99#_c_1627_n N_SLEEP_B_M1020_g 8.27818e-19 $X=15.83 $Y=0.88
+ $X2=0 $Y2=0
cc_1209 N_A_2216_99#_c_1628_n N_SLEEP_B_M1020_g 0.0160934f $X=16.455 $Y=0.965
+ $X2=0 $Y2=0
cc_1210 N_A_2216_99#_c_1630_n N_SLEEP_B_M1020_g 0.0047667f $X=16.645 $Y=1.05
+ $X2=0 $Y2=0
cc_1211 N_A_2216_99#_c_1631_n N_SLEEP_B_M1020_g 0.00136357f $X=16.67 $Y=2.065
+ $X2=0 $Y2=0
cc_1212 N_A_2216_99#_c_1630_n N_SLEEP_B_M1022_g 0.0160999f $X=16.645 $Y=1.05
+ $X2=0 $Y2=0
cc_1213 N_A_2216_99#_c_1631_n N_SLEEP_B_M1022_g 0.00150488f $X=16.67 $Y=2.065
+ $X2=0 $Y2=0
cc_1214 N_A_2216_99#_c_1631_n N_SLEEP_B_c_2167_n 0.00682036f $X=16.67 $Y=2.065
+ $X2=0 $Y2=0
cc_1215 N_A_2216_99#_c_1628_n N_SLEEP_B_c_2168_n 0.0254623f $X=16.455 $Y=0.965
+ $X2=0 $Y2=0
cc_1216 N_A_2216_99#_c_1631_n N_SLEEP_B_c_2168_n 0.0568199f $X=16.67 $Y=2.065
+ $X2=0 $Y2=0
cc_1217 N_A_2216_99#_c_1628_n N_SLEEP_B_c_2169_n 0.00703037f $X=16.455 $Y=0.965
+ $X2=0 $Y2=0
cc_1218 N_A_2216_99#_c_1629_n N_SLEEP_B_c_2169_n 0.0123643f $X=15.915 $Y=0.965
+ $X2=0 $Y2=0
cc_1219 N_A_2216_99#_c_1631_n N_SLEEP_B_c_2169_n 0.031435f $X=16.67 $Y=2.065
+ $X2=0 $Y2=0
cc_1220 N_A_2216_99#_c_1630_n N_A_3466_403#_c_2239_n 0.0130477f $X=16.645
+ $Y=1.05 $X2=0 $Y2=0
cc_1221 N_A_2216_99#_c_1631_n N_A_3466_403#_c_2239_n 0.00407391f $X=16.67
+ $Y=2.065 $X2=0 $Y2=0
cc_1222 N_A_2216_99#_c_1630_n N_A_3466_403#_c_2242_n 0.0191901f $X=16.645
+ $Y=1.05 $X2=0 $Y2=0
cc_1223 N_A_2216_99#_c_1631_n N_A_3466_403#_c_2244_n 0.0104787f $X=16.67
+ $Y=2.065 $X2=0 $Y2=0
cc_1224 N_A_2216_99#_M1024_g N_VPWR_c_2365_n 0.00569155f $X=13.165 $Y=2.57 $X2=0
+ $Y2=0
cc_1225 N_A_2216_99#_M1024_g N_VPWR_c_2354_n 0.00737832f $X=13.165 $Y=2.57 $X2=0
+ $Y2=0
cc_1226 N_A_2216_99#_M1024_g N_KAPWR_c_2675_n 0.0119793f $X=13.165 $Y=2.57 $X2=0
+ $Y2=0
cc_1227 N_A_2216_99#_M1045_d N_KAPWR_c_2677_n 0.00329858f $X=16.53 $Y=1.92 $X2=0
+ $Y2=0
cc_1228 N_A_2216_99#_M1024_g N_KAPWR_c_2677_n 0.00244127f $X=13.165 $Y=2.57
+ $X2=0 $Y2=0
cc_1229 N_A_2216_99#_c_1616_n N_VGND_c_2838_n 0.00305522f $X=11.155 $Y=1.155
+ $X2=0 $Y2=0
cc_1230 N_A_2216_99#_c_1616_n N_VGND_c_2840_n 0.00355641f $X=11.155 $Y=1.155
+ $X2=0 $Y2=0
cc_1231 N_A_2216_99#_c_1621_n N_VGND_c_2840_n 0.0202958f $X=12.165 $Y=1.25 $X2=0
+ $Y2=0
cc_1232 N_A_2216_99#_c_1622_n N_VGND_c_2840_n 0.00486879f $X=11.79 $Y=1.29 $X2=0
+ $Y2=0
cc_1233 N_A_2216_99#_c_1623_n N_VGND_c_2840_n 0.0387097f $X=12.25 $Y=1.125 $X2=0
+ $Y2=0
cc_1234 N_A_2216_99#_c_1625_n N_VGND_c_2840_n 0.0147459f $X=12.335 $Y=0.34 $X2=0
+ $Y2=0
cc_1235 N_A_2216_99#_c_1626_n N_VGND_c_2841_n 0.0113274f $X=15.745 $Y=0.34 $X2=0
+ $Y2=0
cc_1236 N_A_2216_99#_c_1628_n N_VGND_c_2841_n 0.0177054f $X=16.455 $Y=0.965
+ $X2=0 $Y2=0
cc_1237 N_A_2216_99#_c_1630_n N_VGND_c_2841_n 0.00689583f $X=16.645 $Y=1.05
+ $X2=0 $Y2=0
cc_1238 N_A_2216_99#_c_1624_n N_VGND_c_2847_n 0.0766028f $X=13.525 $Y=0.34 $X2=0
+ $Y2=0
cc_1239 N_A_2216_99#_c_1625_n N_VGND_c_2847_n 0.0115893f $X=12.335 $Y=0.34 $X2=0
+ $Y2=0
cc_1240 N_A_2216_99#_c_1626_n N_VGND_c_2847_n 0.132473f $X=15.745 $Y=0.34 $X2=0
+ $Y2=0
cc_1241 N_A_2216_99#_c_1632_n N_VGND_c_2847_n 0.0217908f $X=13.69 $Y=0.34 $X2=0
+ $Y2=0
cc_1242 N_A_2216_99#_c_1630_n N_VGND_c_2852_n 0.012199f $X=16.645 $Y=1.05 $X2=0
+ $Y2=0
cc_1243 N_A_2216_99#_c_1616_n N_VGND_c_2854_n 9.49986e-19 $X=11.155 $Y=1.155
+ $X2=0 $Y2=0
cc_1244 N_A_2216_99#_c_1624_n N_VGND_c_2854_n 0.0399955f $X=13.525 $Y=0.34 $X2=0
+ $Y2=0
cc_1245 N_A_2216_99#_c_1625_n N_VGND_c_2854_n 0.00583135f $X=12.335 $Y=0.34
+ $X2=0 $Y2=0
cc_1246 N_A_2216_99#_c_1626_n N_VGND_c_2854_n 0.0745908f $X=15.745 $Y=0.34 $X2=0
+ $Y2=0
cc_1247 N_A_2216_99#_c_1630_n N_VGND_c_2854_n 0.0146232f $X=16.645 $Y=1.05 $X2=0
+ $Y2=0
cc_1248 N_A_2216_99#_c_1632_n N_VGND_c_2854_n 0.0111356f $X=13.69 $Y=0.34 $X2=0
+ $Y2=0
cc_1249 N_A_2216_99#_c_1616_n N_A_2074_125#_c_3022_n 5.69865e-19 $X=11.155
+ $Y=1.155 $X2=0 $Y2=0
cc_1250 N_A_2216_99#_c_1617_n N_A_2074_125#_c_3023_n 0.0111789f $X=11.23 $Y=1.23
+ $X2=0 $Y2=0
cc_1251 N_A_2216_99#_c_1621_n N_A_2074_125#_c_3023_n 0.0146639f $X=12.165
+ $Y=1.25 $X2=0 $Y2=0
cc_1252 N_A_2216_99#_c_1622_n N_A_2074_125#_c_3023_n 5.46117e-19 $X=11.79
+ $Y=1.29 $X2=0 $Y2=0
cc_1253 N_A_2216_99#_c_1634_n N_A_2074_125#_c_3023_n 0.00543753f $X=11.625
+ $Y=1.29 $X2=0 $Y2=0
cc_1254 N_A_2216_99#_c_1616_n N_A_2074_125#_c_3025_n 0.00978418f $X=11.155
+ $Y=1.155 $X2=0 $Y2=0
cc_1255 N_A_2216_99#_c_1617_n N_A_2074_125#_c_3025_n 9.922e-19 $X=11.23 $Y=1.23
+ $X2=0 $Y2=0
cc_1256 N_A_2216_99#_c_1621_n N_A_2074_125#_c_3025_n 0.00628218f $X=12.165
+ $Y=1.25 $X2=0 $Y2=0
cc_1257 N_A_2216_99#_c_1634_n N_A_2074_125#_c_3025_n 0.00682168f $X=11.625
+ $Y=1.29 $X2=0 $Y2=0
cc_1258 N_A_2216_99#_c_1626_n A_3056_72# 0.00134117f $X=15.745 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1259 N_A_2216_99#_c_1626_n A_3134_72# 6.48644e-19 $X=15.745 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1260 N_A_2216_99#_c_1627_n A_3134_72# 0.00336593f $X=15.83 $Y=0.88 $X2=-0.19
+ $Y2=-0.245
cc_1261 N_A_1728_125#_M1051_g N_SET_B_c_2004_n 0.00974028f $X=12.24 $Y=0.805
+ $X2=0 $Y2=0
cc_1262 N_A_1728_125#_M1041_g N_SET_B_c_2004_n 0.00882199f $X=12.6 $Y=0.805
+ $X2=0 $Y2=0
cc_1263 N_A_1728_125#_c_1830_n N_SET_B_M1043_g 0.0128789f $X=13.8 $Y=2.65 $X2=0
+ $Y2=0
cc_1264 N_A_1728_125#_c_1802_n N_CLK_M1039_g 0.0142521f $X=17.05 $Y=2.405 $X2=0
+ $Y2=0
cc_1265 N_A_1728_125#_c_1802_n CLK 0.0210364f $X=17.05 $Y=2.405 $X2=0 $Y2=0
cc_1266 N_A_1728_125#_c_1802_n N_CLK_c_2123_n 0.00198094f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1267 N_A_1728_125#_c_1802_n N_SLEEP_B_M1026_g 0.0148923f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1268 N_A_1728_125#_c_1802_n N_SLEEP_B_c_2171_n 0.0228399f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1269 N_A_1728_125#_c_1803_n N_SLEEP_B_c_2171_n 0.00337417f $X=17.135 $Y=2.32
+ $X2=0 $Y2=0
cc_1270 N_A_1728_125#_c_1790_n N_SLEEP_B_c_2171_n 9.07704e-19 $X=17.17 $Y=1.66
+ $X2=0 $Y2=0
cc_1271 N_A_1728_125#_c_1786_n N_SLEEP_B_M1022_g 0.00716535f $X=17.335 $Y=0.87
+ $X2=0 $Y2=0
cc_1272 N_A_1728_125#_c_1802_n N_SLEEP_B_c_2168_n 0.0216644f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1273 N_A_1728_125#_c_1784_n N_SLEEP_B_c_2169_n 0.00983879f $X=17.26 $Y=1.495
+ $X2=0 $Y2=0
cc_1274 N_A_1728_125#_c_1789_n N_SLEEP_B_c_2169_n 2.75549e-19 $X=17.17 $Y=1.66
+ $X2=0 $Y2=0
cc_1275 N_A_1728_125#_c_1790_n N_SLEEP_B_c_2169_n 0.0066741f $X=17.17 $Y=1.66
+ $X2=0 $Y2=0
cc_1276 N_A_1728_125#_c_1797_n N_A_3466_403#_M1004_g 0.0159686f $X=17.615
+ $Y=1.83 $X2=0 $Y2=0
cc_1277 N_A_1728_125#_c_1797_n N_A_3466_403#_c_2247_n 0.00507344f $X=17.615
+ $Y=1.83 $X2=0 $Y2=0
cc_1278 N_A_1728_125#_c_1798_n N_A_3466_403#_c_2247_n 0.00218854f $X=17.69
+ $Y=1.905 $X2=0 $Y2=0
cc_1279 N_A_1728_125#_c_1803_n N_A_3466_403#_c_2247_n 0.0249405f $X=17.135
+ $Y=2.32 $X2=0 $Y2=0
cc_1280 N_A_1728_125#_c_1798_n N_A_3466_403#_c_2248_n 0.00792755f $X=17.69
+ $Y=1.905 $X2=0 $Y2=0
cc_1281 N_A_1728_125#_c_1802_n N_A_3466_403#_c_2248_n 0.0146302f $X=17.05
+ $Y=2.405 $X2=0 $Y2=0
cc_1282 N_A_1728_125#_c_1784_n N_A_3466_403#_c_2239_n 0.00359506f $X=17.26
+ $Y=1.495 $X2=0 $Y2=0
cc_1283 N_A_1728_125#_c_1785_n N_A_3466_403#_c_2239_n 0.013693f $X=17.63 $Y=0.87
+ $X2=0 $Y2=0
cc_1284 N_A_1728_125#_M1007_g N_A_3466_403#_c_2239_n 0.00340635f $X=17.705
+ $Y=0.445 $X2=0 $Y2=0
cc_1285 N_A_1728_125#_c_1785_n N_A_3466_403#_c_2240_n 0.00430222f $X=17.63
+ $Y=0.87 $X2=0 $Y2=0
cc_1286 N_A_1728_125#_c_1797_n N_A_3466_403#_c_2240_n 0.00368494f $X=17.615
+ $Y=1.83 $X2=0 $Y2=0
cc_1287 N_A_1728_125#_c_1784_n N_A_3466_403#_c_2241_n 0.0041774f $X=17.26
+ $Y=1.495 $X2=0 $Y2=0
cc_1288 N_A_1728_125#_c_1786_n N_A_3466_403#_c_2242_n 0.00719969f $X=17.335
+ $Y=0.87 $X2=0 $Y2=0
cc_1289 N_A_1728_125#_M1007_g N_A_3466_403#_c_2242_n 0.00570787f $X=17.705
+ $Y=0.445 $X2=0 $Y2=0
cc_1290 N_A_1728_125#_c_1797_n N_A_3466_403#_c_2243_n 0.0130668f $X=17.615
+ $Y=1.83 $X2=0 $Y2=0
cc_1291 N_A_1728_125#_c_1798_n N_A_3466_403#_c_2243_n 0.00258935f $X=17.69
+ $Y=1.905 $X2=0 $Y2=0
cc_1292 N_A_1728_125#_c_1803_n N_A_3466_403#_c_2243_n 0.00827308f $X=17.135
+ $Y=2.32 $X2=0 $Y2=0
cc_1293 N_A_1728_125#_c_1789_n N_A_3466_403#_c_2243_n 0.0230003f $X=17.17
+ $Y=1.66 $X2=0 $Y2=0
cc_1294 N_A_1728_125#_c_1790_n N_A_3466_403#_c_2243_n 0.00336089f $X=17.17
+ $Y=1.66 $X2=0 $Y2=0
cc_1295 N_A_1728_125#_c_1784_n N_A_3466_403#_c_2244_n 0.00521466f $X=17.26
+ $Y=1.495 $X2=0 $Y2=0
cc_1296 N_A_1728_125#_c_1789_n N_A_3466_403#_c_2244_n 0.00168861f $X=17.17
+ $Y=1.66 $X2=0 $Y2=0
cc_1297 N_A_1728_125#_M1007_g N_A_3466_403#_c_2245_n 0.0135565f $X=17.705
+ $Y=0.445 $X2=0 $Y2=0
cc_1298 N_A_1728_125#_c_1797_n N_VPWR_c_2359_n 0.00979444f $X=17.615 $Y=1.83
+ $X2=0 $Y2=0
cc_1299 N_A_1728_125#_c_1795_n N_VPWR_c_2365_n 0.0054269f $X=12.475 $Y=1.895
+ $X2=0 $Y2=0
cc_1300 N_A_1728_125#_c_1798_n N_VPWR_c_2365_n 0.00235582f $X=17.69 $Y=1.905
+ $X2=0 $Y2=0
cc_1301 N_A_1728_125#_c_1823_n N_VPWR_c_2365_n 0.0139169f $X=9.02 $Y=2.62 $X2=0
+ $Y2=0
cc_1302 N_A_1728_125#_c_1801_n N_VPWR_c_2365_n 0.212704f $X=12.315 $Y=2.91 $X2=0
+ $Y2=0
cc_1303 N_A_1728_125#_c_1830_n N_VPWR_c_2365_n 0.00300519f $X=13.8 $Y=2.65 $X2=0
+ $Y2=0
cc_1304 N_A_1728_125#_c_1805_n N_VPWR_c_2365_n 0.0113327f $X=12.4 $Y=2.65 $X2=0
+ $Y2=0
cc_1305 N_A_1728_125#_c_1808_n N_VPWR_c_2365_n 0.00871362f $X=11.3 $Y=2.91 $X2=0
+ $Y2=0
cc_1306 N_A_1728_125#_M1037_d N_VPWR_c_2354_n 0.00121835f $X=8.92 $Y=2.255 $X2=0
+ $Y2=0
cc_1307 N_A_1728_125#_c_1795_n N_VPWR_c_2354_n 0.00661658f $X=12.475 $Y=1.895
+ $X2=0 $Y2=0
cc_1308 N_A_1728_125#_c_1798_n N_VPWR_c_2354_n 7.3165e-19 $X=17.69 $Y=1.905
+ $X2=0 $Y2=0
cc_1309 N_A_1728_125#_c_1823_n N_VPWR_c_2354_n 0.00210636f $X=9.02 $Y=2.62 $X2=0
+ $Y2=0
cc_1310 N_A_1728_125#_c_1801_n N_VPWR_c_2354_n 0.0273741f $X=12.315 $Y=2.91
+ $X2=0 $Y2=0
cc_1311 N_A_1728_125#_c_1830_n N_VPWR_c_2354_n 0.00139559f $X=13.8 $Y=2.65 $X2=0
+ $Y2=0
cc_1312 N_A_1728_125#_c_1805_n N_VPWR_c_2354_n 0.00138619f $X=12.4 $Y=2.65 $X2=0
+ $Y2=0
cc_1313 N_A_1728_125#_c_1808_n N_VPWR_c_2354_n 0.00693807f $X=11.3 $Y=2.91 $X2=0
+ $Y2=0
cc_1314 N_A_1728_125#_c_1830_n N_KAPWR_M1018_d 0.00574979f $X=13.8 $Y=2.65
+ $X2=-0.19 $Y2=-0.245
cc_1315 N_A_1728_125#_c_1802_n N_KAPWR_M1011_d 0.0107789f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1316 N_A_1728_125#_c_1802_n N_KAPWR_M1026_d 0.00595627f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1317 N_A_1728_125#_M1043_d N_KAPWR_c_2675_n 7.82306e-19 $X=13.78 $Y=2.07
+ $X2=0 $Y2=0
cc_1318 N_A_1728_125#_c_1795_n N_KAPWR_c_2675_n 0.00143708f $X=12.475 $Y=1.895
+ $X2=0 $Y2=0
cc_1319 N_A_1728_125#_c_1830_n N_KAPWR_c_2675_n 0.070453f $X=13.8 $Y=2.65 $X2=0
+ $Y2=0
cc_1320 N_A_1728_125#_c_1802_n N_KAPWR_c_2675_n 0.00524821f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1321 N_A_1728_125#_c_1805_n N_KAPWR_c_2675_n 0.0095593f $X=12.4 $Y=2.65 $X2=0
+ $Y2=0
cc_1322 N_A_1728_125#_c_1844_n N_KAPWR_c_2675_n 0.0194814f $X=13.965 $Y=2.435
+ $X2=0 $Y2=0
cc_1323 N_A_1728_125#_c_1847_n N_KAPWR_c_2675_n 0.00880992f $X=14.425 $Y=2.42
+ $X2=0 $Y2=0
cc_1324 N_A_1728_125#_c_1802_n N_KAPWR_c_2676_n 0.0193675f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1325 N_A_1728_125#_M1037_d N_KAPWR_c_2677_n 0.00121402f $X=8.92 $Y=2.255
+ $X2=0 $Y2=0
cc_1326 N_A_1728_125#_c_1791_n N_KAPWR_c_2677_n 0.00356333f $X=11.3 $Y=2.745
+ $X2=0 $Y2=0
cc_1327 N_A_1728_125#_c_1795_n N_KAPWR_c_2677_n 0.0025654f $X=12.475 $Y=1.895
+ $X2=0 $Y2=0
cc_1328 N_A_1728_125#_c_1798_n N_KAPWR_c_2677_n 0.00895912f $X=17.69 $Y=1.905
+ $X2=0 $Y2=0
cc_1329 N_A_1728_125#_c_1823_n N_KAPWR_c_2677_n 0.0223168f $X=9.02 $Y=2.62 $X2=0
+ $Y2=0
cc_1330 N_A_1728_125#_c_1801_n N_KAPWR_c_2677_n 0.11294f $X=12.315 $Y=2.91 $X2=0
+ $Y2=0
cc_1331 N_A_1728_125#_c_1830_n N_KAPWR_c_2677_n 0.0410343f $X=13.8 $Y=2.65 $X2=0
+ $Y2=0
cc_1332 N_A_1728_125#_c_1802_n N_KAPWR_c_2677_n 0.0892003f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1333 N_A_1728_125#_c_1805_n N_KAPWR_c_2677_n 0.0159702f $X=12.4 $Y=2.65 $X2=0
+ $Y2=0
cc_1334 N_A_1728_125#_c_1844_n N_KAPWR_c_2677_n 0.012895f $X=13.965 $Y=2.435
+ $X2=0 $Y2=0
cc_1335 N_A_1728_125#_c_1847_n N_KAPWR_c_2677_n 0.013942f $X=14.425 $Y=2.42
+ $X2=0 $Y2=0
cc_1336 N_A_1728_125#_c_1808_n N_KAPWR_c_2677_n 0.00202167f $X=11.3 $Y=2.91
+ $X2=0 $Y2=0
cc_1337 N_A_1728_125#_c_1802_n N_KAPWR_c_2678_n 0.0235255f $X=17.05 $Y=2.405
+ $X2=0 $Y2=0
cc_1338 N_A_1728_125#_c_1830_n A_2658_414# 0.00252257f $X=13.8 $Y=2.65 $X2=-0.19
+ $Y2=-0.245
cc_1339 N_A_1728_125#_c_1847_n A_2862_414# 0.0028347f $X=14.425 $Y=2.42
+ $X2=-0.19 $Y2=-0.245
cc_1340 N_A_1728_125#_c_1849_n A_2862_414# 0.00553698f $X=14.595 $Y=2.42
+ $X2=-0.19 $Y2=-0.245
cc_1341 N_A_1728_125#_M1051_g N_VGND_c_2840_n 0.00945444f $X=12.24 $Y=0.805
+ $X2=0 $Y2=0
cc_1342 N_A_1728_125#_M1007_g N_VGND_c_2842_n 0.0102962f $X=17.705 $Y=0.445
+ $X2=0 $Y2=0
cc_1343 N_A_1728_125#_M1007_g N_VGND_c_2852_n 0.00521005f $X=17.705 $Y=0.445
+ $X2=0 $Y2=0
cc_1344 N_A_1728_125#_c_1786_n N_VGND_c_2854_n 0.00371149f $X=17.335 $Y=0.87
+ $X2=0 $Y2=0
cc_1345 N_A_1728_125#_M1007_g N_VGND_c_2854_n 0.0109789f $X=17.705 $Y=0.445
+ $X2=0 $Y2=0
cc_1346 N_SET_B_M1027_g N_VPWR_c_2358_n 0.00619142f $X=7.06 $Y=2.465 $X2=0 $Y2=0
cc_1347 N_SET_B_M1027_g N_VPWR_c_2364_n 0.00264846f $X=7.06 $Y=2.465 $X2=0 $Y2=0
cc_1348 N_SET_B_M1043_g N_VPWR_c_2365_n 0.00569155f $X=13.655 $Y=2.57 $X2=0
+ $Y2=0
cc_1349 N_SET_B_M1027_g N_VPWR_c_2354_n 7.49299e-19 $X=7.06 $Y=2.465 $X2=0 $Y2=0
cc_1350 N_SET_B_M1043_g N_VPWR_c_2354_n 0.00660084f $X=13.655 $Y=2.57 $X2=0
+ $Y2=0
cc_1351 N_SET_B_M1043_g N_KAPWR_c_2675_n 0.0114841f $X=13.655 $Y=2.57 $X2=0
+ $Y2=0
cc_1352 N_SET_B_M1027_g N_KAPWR_c_2677_n 0.00573698f $X=7.06 $Y=2.465 $X2=0
+ $Y2=0
cc_1353 N_SET_B_M1043_g N_KAPWR_c_2677_n 0.00200246f $X=13.655 $Y=2.57 $X2=0
+ $Y2=0
cc_1354 N_SET_B_M1003_g N_VGND_c_2837_n 0.00895129f $X=7 $Y=0.695 $X2=0 $Y2=0
cc_1355 N_SET_B_c_2001_n N_VGND_c_2837_n 0.0198212f $X=10.65 $Y=0.18 $X2=0 $Y2=0
cc_1356 N_SET_B_M1008_g N_VGND_c_2838_n 0.0170303f $X=10.725 $Y=0.835 $X2=0
+ $Y2=0
cc_1357 N_SET_B_c_2004_n N_VGND_c_2838_n 0.0142544f $X=14.065 $Y=0.18 $X2=0
+ $Y2=0
cc_1358 N_SET_B_c_2009_n N_VGND_c_2838_n 0.00459621f $X=10.725 $Y=0.18 $X2=0
+ $Y2=0
cc_1359 N_SET_B_c_2004_n N_VGND_c_2839_n 0.0226526f $X=14.065 $Y=0.18 $X2=0
+ $Y2=0
cc_1360 N_SET_B_c_2004_n N_VGND_c_2840_n 0.0215559f $X=14.065 $Y=0.18 $X2=0
+ $Y2=0
cc_1361 N_SET_B_c_2002_n N_VGND_c_2845_n 0.00737585f $X=7.075 $Y=0.18 $X2=0
+ $Y2=0
cc_1362 N_SET_B_c_2004_n N_VGND_c_2847_n 0.0481494f $X=14.065 $Y=0.18 $X2=0
+ $Y2=0
cc_1363 N_SET_B_c_2001_n N_VGND_c_2851_n 0.0780065f $X=10.65 $Y=0.18 $X2=0 $Y2=0
cc_1364 N_SET_B_c_2001_n N_VGND_c_2854_n 0.0894887f $X=10.65 $Y=0.18 $X2=0 $Y2=0
cc_1365 N_SET_B_c_2002_n N_VGND_c_2854_n 0.0114428f $X=7.075 $Y=0.18 $X2=0 $Y2=0
cc_1366 N_SET_B_c_2004_n N_VGND_c_2854_n 0.088517f $X=14.065 $Y=0.18 $X2=0 $Y2=0
cc_1367 N_SET_B_c_2009_n N_VGND_c_2854_n 0.00749832f $X=10.725 $Y=0.18 $X2=0
+ $Y2=0
cc_1368 N_SET_B_c_2001_n N_A_2074_125#_c_3022_n 0.00265981f $X=10.65 $Y=0.18
+ $X2=0 $Y2=0
cc_1369 N_SET_B_M1008_g N_A_2074_125#_c_3022_n 0.00187455f $X=10.725 $Y=0.835
+ $X2=0 $Y2=0
cc_1370 N_SET_B_M1008_g N_A_2074_125#_c_3023_n 0.00347642f $X=10.725 $Y=0.835
+ $X2=0 $Y2=0
cc_1371 N_SET_B_M1008_g N_A_2074_125#_c_3025_n 5.72994e-19 $X=10.725 $Y=0.835
+ $X2=0 $Y2=0
cc_1372 N_SET_B_c_2004_n N_A_2074_125#_c_3025_n 0.00451709f $X=14.065 $Y=0.18
+ $X2=0 $Y2=0
cc_1373 N_CLK_M1015_g N_SLEEP_B_M1014_g 0.0464943f $X=15.205 $Y=0.57 $X2=0 $Y2=0
cc_1374 N_CLK_c_2123_n N_SLEEP_B_M1026_g 0.0358292f $X=15.385 $Y=1.51 $X2=0
+ $Y2=0
cc_1375 N_CLK_M1015_g N_SLEEP_B_c_2169_n 0.00587992f $X=15.205 $Y=0.57 $X2=0
+ $Y2=0
cc_1376 N_CLK_c_2123_n N_SLEEP_B_c_2169_n 0.0134798f $X=15.385 $Y=1.51 $X2=0
+ $Y2=0
cc_1377 N_CLK_M1039_g N_VPWR_c_2365_n 0.00228063f $X=15.385 $Y=2.24 $X2=0 $Y2=0
cc_1378 N_CLK_M1039_g N_VPWR_c_2354_n 6.56441e-19 $X=15.385 $Y=2.24 $X2=0 $Y2=0
cc_1379 CLK N_KAPWR_M1011_d 0.0108074f $X=15.035 $Y=1.21 $X2=0 $Y2=0
cc_1380 N_CLK_M1039_g N_KAPWR_c_2677_n 0.00356477f $X=15.385 $Y=2.24 $X2=0 $Y2=0
cc_1381 N_CLK_M1039_g N_KAPWR_c_2678_n 7.75614e-19 $X=15.385 $Y=2.24 $X2=0 $Y2=0
cc_1382 N_CLK_M1015_g N_VGND_c_2847_n 0.00283474f $X=15.205 $Y=0.57 $X2=0 $Y2=0
cc_1383 N_CLK_M1015_g N_VGND_c_2854_n 0.00385656f $X=15.205 $Y=0.57 $X2=0 $Y2=0
cc_1384 N_SLEEP_B_M1022_g N_A_3466_403#_c_2239_n 7.35457e-19 $X=16.745 $Y=0.57
+ $X2=0 $Y2=0
cc_1385 N_SLEEP_B_M1022_g N_A_3466_403#_c_2242_n 0.00275298f $X=16.745 $Y=0.57
+ $X2=0 $Y2=0
cc_1386 N_SLEEP_B_M1026_g N_VPWR_c_2365_n 0.00228063f $X=15.815 $Y=2.24 $X2=0
+ $Y2=0
cc_1387 N_SLEEP_B_c_2171_n N_VPWR_c_2365_n 0.00888725f $X=16.405 $Y=1.915 $X2=0
+ $Y2=0
cc_1388 N_SLEEP_B_M1026_g N_VPWR_c_2354_n 6.56441e-19 $X=15.815 $Y=2.24 $X2=0
+ $Y2=0
cc_1389 N_SLEEP_B_c_2171_n N_VPWR_c_2354_n 0.00520432f $X=16.405 $Y=1.915 $X2=0
+ $Y2=0
cc_1390 N_SLEEP_B_c_2168_n N_KAPWR_M1026_d 0.00639218f $X=16.095 $Y=1.385 $X2=0
+ $Y2=0
cc_1391 N_SLEEP_B_M1026_g N_KAPWR_c_2676_n 7.24911e-19 $X=15.815 $Y=2.24 $X2=0
+ $Y2=0
cc_1392 N_SLEEP_B_c_2171_n N_KAPWR_c_2676_n 0.00756886f $X=16.405 $Y=1.915 $X2=0
+ $Y2=0
cc_1393 N_SLEEP_B_M1026_g N_KAPWR_c_2677_n 0.00354408f $X=15.815 $Y=2.24 $X2=0
+ $Y2=0
cc_1394 N_SLEEP_B_c_2171_n N_KAPWR_c_2677_n 0.00896402f $X=16.405 $Y=1.915 $X2=0
+ $Y2=0
cc_1395 N_SLEEP_B_M1049_g N_VGND_c_2841_n 0.00133018f $X=15.955 $Y=0.57 $X2=0
+ $Y2=0
cc_1396 N_SLEEP_B_M1020_g N_VGND_c_2841_n 0.00967933f $X=16.385 $Y=0.57 $X2=0
+ $Y2=0
cc_1397 N_SLEEP_B_M1022_g N_VGND_c_2841_n 0.00166273f $X=16.745 $Y=0.57 $X2=0
+ $Y2=0
cc_1398 N_SLEEP_B_M1014_g N_VGND_c_2847_n 0.00283474f $X=15.595 $Y=0.57 $X2=0
+ $Y2=0
cc_1399 N_SLEEP_B_M1049_g N_VGND_c_2847_n 0.00426187f $X=15.955 $Y=0.57 $X2=0
+ $Y2=0
cc_1400 N_SLEEP_B_M1020_g N_VGND_c_2852_n 0.00389963f $X=16.385 $Y=0.57 $X2=0
+ $Y2=0
cc_1401 N_SLEEP_B_M1022_g N_VGND_c_2852_n 0.00327705f $X=16.745 $Y=0.57 $X2=0
+ $Y2=0
cc_1402 N_SLEEP_B_M1014_g N_VGND_c_2854_n 0.00368401f $X=15.595 $Y=0.57 $X2=0
+ $Y2=0
cc_1403 N_SLEEP_B_M1049_g N_VGND_c_2854_n 0.00792494f $X=15.955 $Y=0.57 $X2=0
+ $Y2=0
cc_1404 N_SLEEP_B_M1020_g N_VGND_c_2854_n 0.00762433f $X=16.385 $Y=0.57 $X2=0
+ $Y2=0
cc_1405 N_SLEEP_B_M1022_g N_VGND_c_2854_n 0.00435779f $X=16.745 $Y=0.57 $X2=0
+ $Y2=0
cc_1406 N_A_3466_403#_M1004_g N_VPWR_c_2359_n 0.0223763f $X=18.235 $Y=2.465
+ $X2=0 $Y2=0
cc_1407 N_A_3466_403#_c_2240_n N_VPWR_c_2359_n 0.0183335f $X=18.095 $Y=1.35
+ $X2=0 $Y2=0
cc_1408 N_A_3466_403#_c_2241_n N_VPWR_c_2359_n 0.00497129f $X=18.095 $Y=1.35
+ $X2=0 $Y2=0
cc_1409 N_A_3466_403#_c_2243_n N_VPWR_c_2359_n 0.0629471f $X=17.532 $Y=1.995
+ $X2=0 $Y2=0
cc_1410 N_A_3466_403#_c_2248_n N_VPWR_c_2365_n 0.00517105f $X=17.475 $Y=2.16
+ $X2=0 $Y2=0
cc_1411 N_A_3466_403#_M1004_g N_VPWR_c_2366_n 0.00486043f $X=18.235 $Y=2.465
+ $X2=0 $Y2=0
cc_1412 N_A_3466_403#_M1004_g N_VPWR_c_2354_n 0.00453305f $X=18.235 $Y=2.465
+ $X2=0 $Y2=0
cc_1413 N_A_3466_403#_c_2248_n N_VPWR_c_2354_n 9.0945e-19 $X=17.475 $Y=2.16
+ $X2=0 $Y2=0
cc_1414 N_A_3466_403#_M1004_g N_KAPWR_c_2677_n 0.00675489f $X=18.235 $Y=2.465
+ $X2=0 $Y2=0
cc_1415 N_A_3466_403#_c_2248_n N_KAPWR_c_2677_n 0.0127266f $X=17.475 $Y=2.16
+ $X2=0 $Y2=0
cc_1416 N_A_3466_403#_M1004_g N_Q_c_2818_n 0.0157653f $X=18.235 $Y=2.465 $X2=0
+ $Y2=0
cc_1417 N_A_3466_403#_c_2240_n N_Q_c_2818_n 0.0270266f $X=18.095 $Y=1.35 $X2=0
+ $Y2=0
cc_1418 N_A_3466_403#_c_2245_n N_Q_c_2818_n 0.0157061f $X=18.122 $Y=1.185 $X2=0
+ $Y2=0
cc_1419 N_A_3466_403#_c_2240_n N_VGND_c_2842_n 0.024755f $X=18.095 $Y=1.35 $X2=0
+ $Y2=0
cc_1420 N_A_3466_403#_c_2241_n N_VGND_c_2842_n 0.00532052f $X=18.095 $Y=1.35
+ $X2=0 $Y2=0
cc_1421 N_A_3466_403#_c_2242_n N_VGND_c_2842_n 0.0520862f $X=17.49 $Y=0.445
+ $X2=0 $Y2=0
cc_1422 N_A_3466_403#_c_2245_n N_VGND_c_2842_n 0.0150721f $X=18.122 $Y=1.185
+ $X2=0 $Y2=0
cc_1423 N_A_3466_403#_c_2242_n N_VGND_c_2852_n 0.0174241f $X=17.49 $Y=0.445
+ $X2=0 $Y2=0
cc_1424 N_A_3466_403#_c_2245_n N_VGND_c_2853_n 0.00486043f $X=18.122 $Y=1.185
+ $X2=0 $Y2=0
cc_1425 N_A_3466_403#_M1007_s N_VGND_c_2854_n 0.00222165f $X=17.36 $Y=0.235
+ $X2=0 $Y2=0
cc_1426 N_A_3466_403#_c_2242_n N_VGND_c_2854_n 0.0129307f $X=17.49 $Y=0.445
+ $X2=0 $Y2=0
cc_1427 N_A_3466_403#_c_2245_n N_VGND_c_2854_n 0.00918457f $X=18.122 $Y=1.185
+ $X2=0 $Y2=0
cc_1428 N_A_27_481#_c_2300_n N_VPWR_c_2355_n 0.030529f $X=0.265 $Y=2.55 $X2=0
+ $Y2=0
cc_1429 N_A_27_481#_c_2301_n N_VPWR_c_2355_n 0.0198997f $X=1.02 $Y=2.13 $X2=0
+ $Y2=0
cc_1430 N_A_27_481#_c_2303_n N_VPWR_c_2355_n 0.0364226f $X=1.105 $Y=2.905 $X2=0
+ $Y2=0
cc_1431 N_A_27_481#_c_2305_n N_VPWR_c_2355_n 0.01326f $X=1.19 $Y=2.99 $X2=0
+ $Y2=0
cc_1432 N_A_27_481#_c_2300_n N_VPWR_c_2362_n 0.0220321f $X=0.265 $Y=2.55 $X2=0
+ $Y2=0
cc_1433 N_A_27_481#_c_2304_n N_VPWR_c_2363_n 0.0649237f $X=1.94 $Y=2.99 $X2=0
+ $Y2=0
cc_1434 N_A_27_481#_c_2305_n N_VPWR_c_2363_n 0.0119959f $X=1.19 $Y=2.99 $X2=0
+ $Y2=0
cc_1435 N_A_27_481#_c_2300_n N_VPWR_c_2354_n 0.0030822f $X=0.265 $Y=2.55 $X2=0
+ $Y2=0
cc_1436 N_A_27_481#_c_2304_n N_VPWR_c_2354_n 0.00806174f $X=1.94 $Y=2.99 $X2=0
+ $Y2=0
cc_1437 N_A_27_481#_c_2305_n N_VPWR_c_2354_n 0.00154424f $X=1.19 $Y=2.99 $X2=0
+ $Y2=0
cc_1438 N_A_27_481#_c_2303_n A_213_481# 0.00581947f $X=1.105 $Y=2.905 $X2=-0.19
+ $Y2=1.655
cc_1439 N_A_27_481#_c_2304_n A_213_481# 9.71172e-19 $X=1.94 $Y=2.99 $X2=-0.19
+ $Y2=1.655
cc_1440 N_A_27_481#_c_2304_n N_A_189_119#_M1012_d 7.82306e-19 $X=1.94 $Y=2.99
+ $X2=0 $Y2=0
cc_1441 N_A_27_481#_c_2304_n N_A_189_119#_c_2526_n 0.00237888f $X=1.94 $Y=2.99
+ $X2=0 $Y2=0
cc_1442 N_A_27_481#_c_2306_n N_A_189_119#_c_2526_n 0.0187091f $X=2.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1443 N_A_27_481#_c_2303_n N_A_189_119#_c_2531_n 0.0285796f $X=1.105 $Y=2.905
+ $X2=0 $Y2=0
cc_1444 N_A_27_481#_c_2304_n N_A_189_119#_c_2531_n 0.0196167f $X=1.94 $Y=2.99
+ $X2=0 $Y2=0
cc_1445 N_A_27_481#_c_2306_n N_A_189_119#_c_2531_n 0.00717549f $X=2.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1446 N_A_27_481#_c_2301_n N_A_189_119#_c_2525_n 0.00775699f $X=1.02 $Y=2.13
+ $X2=0 $Y2=0
cc_1447 N_A_27_481#_c_2303_n N_A_189_119#_c_2525_n 3.6704e-19 $X=1.105 $Y=2.905
+ $X2=0 $Y2=0
cc_1448 N_A_27_481#_M1048_d N_KAPWR_c_2677_n 5.07094e-19 $X=1.885 $Y=2.405 $X2=0
+ $Y2=0
cc_1449 N_A_27_481#_c_2300_n N_KAPWR_c_2677_n 0.0387481f $X=0.265 $Y=2.55 $X2=0
+ $Y2=0
cc_1450 N_A_27_481#_c_2301_n N_KAPWR_c_2677_n 0.011525f $X=1.02 $Y=2.13 $X2=0
+ $Y2=0
cc_1451 N_A_27_481#_c_2303_n N_KAPWR_c_2677_n 0.0218782f $X=1.105 $Y=2.905 $X2=0
+ $Y2=0
cc_1452 N_A_27_481#_c_2304_n N_KAPWR_c_2677_n 0.0252256f $X=1.94 $Y=2.99 $X2=0
+ $Y2=0
cc_1453 N_A_27_481#_c_2305_n N_KAPWR_c_2677_n 0.00249508f $X=1.19 $Y=2.99 $X2=0
+ $Y2=0
cc_1454 N_A_27_481#_c_2306_n N_KAPWR_c_2677_n 0.0239236f $X=2.025 $Y=2.815 $X2=0
+ $Y2=0
cc_1455 N_VPWR_c_2354_n N_A_189_119#_M1005_s 0.00168871f $X=18.48 $Y=3.33 $X2=0
+ $Y2=0
cc_1456 N_VPWR_M1036_d N_A_189_119#_c_2526_n 0.0190202f $X=2.845 $Y=1.795 $X2=0
+ $Y2=0
cc_1457 N_VPWR_c_2356_n N_A_189_119#_c_2526_n 0.0250875f $X=3.085 $Y=2.73 $X2=0
+ $Y2=0
cc_1458 N_VPWR_c_2356_n N_A_189_119#_c_2527_n 0.00381204f $X=3.085 $Y=2.73 $X2=0
+ $Y2=0
cc_1459 N_VPWR_c_2360_n N_A_189_119#_c_2528_n 0.0165623f $X=6.025 $Y=3.33 $X2=0
+ $Y2=0
cc_1460 N_VPWR_c_2354_n N_A_189_119#_c_2528_n 0.00205919f $X=18.48 $Y=3.33 $X2=0
+ $Y2=0
cc_1461 N_VPWR_c_2356_n N_A_189_119#_c_2529_n 0.00534229f $X=3.085 $Y=2.73 $X2=0
+ $Y2=0
cc_1462 N_VPWR_c_2360_n N_A_189_119#_c_2529_n 0.00484993f $X=6.025 $Y=3.33 $X2=0
+ $Y2=0
cc_1463 N_VPWR_c_2354_n N_A_189_119#_c_2529_n 5.75857e-19 $X=18.48 $Y=3.33 $X2=0
+ $Y2=0
cc_1464 N_VPWR_c_2360_n N_A_189_119#_c_2523_n 0.0341672f $X=6.025 $Y=3.33 $X2=0
+ $Y2=0
cc_1465 N_VPWR_c_2354_n N_A_189_119#_c_2523_n 0.00445671f $X=18.48 $Y=3.33 $X2=0
+ $Y2=0
cc_1466 N_VPWR_c_2354_n A_1132_535# 0.00194712f $X=18.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1467 N_VPWR_c_2354_n N_A_1541_125#_M1032_d 0.00319411f $X=18.48 $Y=3.33 $X2=0
+ $Y2=0
cc_1468 N_VPWR_c_2354_n A_1712_451# 0.00115927f $X=18.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1469 N_VPWR_c_2354_n N_KAPWR_M1018_d 0.00131774f $X=18.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1470 N_VPWR_c_2365_n N_KAPWR_c_2675_n 0.141731f $X=17.855 $Y=3.33 $X2=0 $Y2=0
cc_1471 N_VPWR_c_2354_n N_KAPWR_c_2675_n 0.0172702f $X=18.48 $Y=3.33 $X2=0 $Y2=0
cc_1472 N_VPWR_c_2365_n N_KAPWR_c_2676_n 0.0134999f $X=17.855 $Y=3.33 $X2=0
+ $Y2=0
cc_1473 N_VPWR_c_2354_n N_KAPWR_c_2676_n 0.0014932f $X=18.48 $Y=3.33 $X2=0 $Y2=0
cc_1474 N_VPWR_M1000_d N_KAPWR_c_2677_n 0.00183293f $X=0.555 $Y=2.405 $X2=0
+ $Y2=0
cc_1475 N_VPWR_M1035_d N_KAPWR_c_2677_n 0.00115506f $X=6.05 $Y=2.675 $X2=0 $Y2=0
cc_1476 N_VPWR_M1027_d N_KAPWR_c_2677_n 0.00158417f $X=7.135 $Y=2.255 $X2=0
+ $Y2=0
cc_1477 N_VPWR_c_2355_n N_KAPWR_c_2677_n 0.0204245f $X=0.765 $Y=2.55 $X2=0 $Y2=0
cc_1478 N_VPWR_c_2356_n N_KAPWR_c_2677_n 0.0350612f $X=3.085 $Y=2.73 $X2=0 $Y2=0
cc_1479 N_VPWR_c_2357_n N_KAPWR_c_2677_n 0.0316853f $X=6.19 $Y=2.885 $X2=0 $Y2=0
cc_1480 N_VPWR_c_2358_n N_KAPWR_c_2677_n 0.0333902f $X=7.415 $Y=2.42 $X2=0 $Y2=0
cc_1481 N_VPWR_c_2359_n N_KAPWR_c_2677_n 0.0447483f $X=18.02 $Y=1.98 $X2=0 $Y2=0
cc_1482 N_VPWR_c_2360_n N_KAPWR_c_2677_n 0.0088807f $X=6.025 $Y=3.33 $X2=0 $Y2=0
cc_1483 N_VPWR_c_2362_n N_KAPWR_c_2677_n 0.00126129f $X=0.6 $Y=3.33 $X2=0 $Y2=0
cc_1484 N_VPWR_c_2363_n N_KAPWR_c_2677_n 0.00557094f $X=2.92 $Y=3.33 $X2=0 $Y2=0
cc_1485 N_VPWR_c_2364_n N_KAPWR_c_2677_n 0.0040129f $X=7.25 $Y=3.33 $X2=0 $Y2=0
cc_1486 N_VPWR_c_2365_n N_KAPWR_c_2677_n 0.0197147f $X=17.855 $Y=3.33 $X2=0
+ $Y2=0
cc_1487 N_VPWR_c_2366_n N_KAPWR_c_2677_n 0.00125273f $X=18.48 $Y=3.33 $X2=0
+ $Y2=0
cc_1488 N_VPWR_c_2354_n N_KAPWR_c_2677_n 1.95712f $X=18.48 $Y=3.33 $X2=0 $Y2=0
cc_1489 N_VPWR_c_2365_n N_KAPWR_c_2678_n 0.0226635f $X=17.855 $Y=3.33 $X2=0
+ $Y2=0
cc_1490 N_VPWR_c_2354_n N_KAPWR_c_2678_n 0.00292358f $X=18.48 $Y=3.33 $X2=0
+ $Y2=0
cc_1491 N_VPWR_c_2354_n N_Q_M1004_d 0.00137166f $X=18.48 $Y=3.33 $X2=0 $Y2=0
cc_1492 N_VPWR_c_2359_n N_Q_c_2818_n 0.0490351f $X=18.02 $Y=1.98 $X2=0 $Y2=0
cc_1493 N_VPWR_c_2366_n N_Q_c_2818_n 0.017801f $X=18.48 $Y=3.33 $X2=0 $Y2=0
cc_1494 N_VPWR_c_2354_n N_Q_c_2818_n 0.00237217f $X=18.48 $Y=3.33 $X2=0 $Y2=0
cc_1495 A_213_481# N_KAPWR_c_2677_n 0.00469538f $X=1.065 $Y=2.405 $X2=2.065
+ $Y2=2.815
cc_1496 N_A_189_119#_M1005_s N_KAPWR_c_2677_n 8.28993e-19 $X=4.725 $Y=2.675
+ $X2=0 $Y2=0
cc_1497 N_A_189_119#_c_2526_n N_KAPWR_c_2677_n 0.0558109f $X=3.665 $Y=2.31 $X2=0
+ $Y2=0
cc_1498 N_A_189_119#_c_2528_n N_KAPWR_c_2677_n 0.0314137f $X=4.43 $Y=2.74 $X2=0
+ $Y2=0
cc_1499 N_A_189_119#_c_2529_n N_KAPWR_c_2677_n 0.0165339f $X=3.835 $Y=2.74 $X2=0
+ $Y2=0
cc_1500 N_A_189_119#_c_2523_n N_KAPWR_c_2677_n 0.0419088f $X=4.515 $Y=2.655
+ $X2=0 $Y2=0
cc_1501 N_A_189_119#_c_2531_n N_KAPWR_c_2677_n 0.0249569f $X=1.6 $Y=2.31 $X2=0
+ $Y2=0
cc_1502 N_A_189_119#_c_2524_n N_VGND_c_2833_n 0.0145731f $X=1.085 $Y=0.805 $X2=0
+ $Y2=0
cc_1503 N_A_189_119#_c_2519_n N_VGND_c_2834_n 0.0134758f $X=1.6 $Y=0.95 $X2=0
+ $Y2=0
cc_1504 N_A_189_119#_c_2524_n N_VGND_c_2843_n 0.00723201f $X=1.085 $Y=0.805
+ $X2=0 $Y2=0
cc_1505 N_A_189_119#_c_2519_n N_VGND_c_2854_n 0.0056259f $X=1.6 $Y=0.95 $X2=0
+ $Y2=0
cc_1506 N_A_189_119#_c_2524_n N_VGND_c_2854_n 0.0088491f $X=1.085 $Y=0.805 $X2=0
+ $Y2=0
cc_1507 N_A_189_119#_c_2519_n A_275_119# 0.0032305f $X=1.6 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_1508 A_1132_535# N_KAPWR_c_2677_n 0.00452178f $X=5.66 $Y=2.675 $X2=0.765
+ $Y2=2.55
cc_1509 N_A_1541_125#_M1032_d N_KAPWR_c_2677_n 0.0170218f $X=7.705 $Y=2.255
+ $X2=0 $Y2=0
cc_1510 N_A_1541_125#_c_2637_n N_KAPWR_c_2677_n 0.00586714f $X=8.27 $Y=2.4 $X2=0
+ $Y2=0
cc_1511 N_A_1541_125#_c_2653_n A_1656_125# 0.00185401f $X=8.27 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_1512 A_1712_451# N_KAPWR_c_2677_n 0.00344388f $X=8.56 $Y=2.255 $X2=8.205
+ $Y2=1.41
cc_1513 N_KAPWR_c_2675_n A_2658_414# 5.92614e-19 $X=14.905 $Y=2.99 $X2=-0.19
+ $Y2=1.655
cc_1514 N_KAPWR_c_2675_n A_2862_414# 0.00148845f $X=14.905 $Y=2.99 $X2=-0.19
+ $Y2=1.655
cc_1515 N_KAPWR_c_2677_n A_2862_414# 0.00223429f $X=16.08 $Y=2.82 $X2=-0.19
+ $Y2=1.655
cc_1516 N_KAPWR_c_2677_n N_Q_M1004_d 0.00244555f $X=16.08 $Y=2.82 $X2=0 $Y2=0
cc_1517 N_KAPWR_c_2677_n N_Q_c_2818_n 0.0320927f $X=16.08 $Y=2.82 $X2=0 $Y2=0
cc_1518 N_Q_c_2818_n N_VGND_c_2853_n 0.0176268f $X=18.455 $Y=0.42 $X2=0 $Y2=0
cc_1519 N_Q_M1033_d N_VGND_c_2854_n 0.00393285f $X=18.315 $Y=0.235 $X2=0 $Y2=0
cc_1520 N_Q_c_2818_n N_VGND_c_2854_n 0.00983606f $X=18.455 $Y=0.42 $X2=0 $Y2=0
cc_1521 N_VGND_c_2854_n A_996_73# 0.00409769f $X=18.48 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1522 N_VGND_c_2838_n N_A_2074_125#_c_3022_n 0.0154564f $X=10.94 $Y=0.82 $X2=0
+ $Y2=0
cc_1523 N_VGND_c_2851_n N_A_2074_125#_c_3022_n 0.0036205f $X=10.775 $Y=0 $X2=0
+ $Y2=0
cc_1524 N_VGND_c_2854_n N_A_2074_125#_c_3022_n 0.0045483f $X=18.48 $Y=0 $X2=0
+ $Y2=0
cc_1525 N_VGND_c_2838_n N_A_2074_125#_c_3023_n 0.017837f $X=10.94 $Y=0.82 $X2=0
+ $Y2=0
cc_1526 N_VGND_c_2838_n N_A_2074_125#_c_3025_n 0.0154978f $X=10.94 $Y=0.82 $X2=0
+ $Y2=0
cc_1527 N_VGND_c_2839_n N_A_2074_125#_c_3025_n 0.00528689f $X=11.745 $Y=0 $X2=0
+ $Y2=0
cc_1528 N_VGND_c_2840_n N_A_2074_125#_c_3025_n 0.0187688f $X=11.91 $Y=0.765
+ $X2=0 $Y2=0
cc_1529 N_VGND_c_2854_n N_A_2074_125#_c_3025_n 0.00668574f $X=18.48 $Y=0 $X2=0
+ $Y2=0
