# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a41oi_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a41oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065000 1.405000 4.095000 1.575000 ;
        RECT 2.555000 1.210000 3.205000 1.405000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.625000 1.195000 5.975000 1.585000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.185000 1.315000 7.535000 1.355000 ;
        RECT 6.185000 1.355000 8.215000 1.585000 ;
        RECT 7.345000 1.155000 7.535000 1.315000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.425000 1.200000 10.455000 1.585000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.210000 1.825000 1.435000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.605000 1.815000 1.745000 ;
        RECT 0.540000 1.745000 4.455000 1.790000 ;
        RECT 0.540000 1.790000 0.870000 2.735000 ;
        RECT 0.595000 0.255000 0.785000 0.855000 ;
        RECT 0.595000 0.855000 3.970000 1.040000 ;
        RECT 1.400000 1.790000 4.455000 1.935000 ;
        RECT 1.400000 1.935000 1.730000 2.735000 ;
        RECT 1.455000 0.255000 1.645000 0.815000 ;
        RECT 1.455000 0.815000 3.970000 0.855000 ;
        RECT 3.640000 0.595000 3.970000 0.815000 ;
        RECT 3.640000 1.040000 3.970000 1.065000 ;
        RECT 3.640000 1.065000 4.455000 1.235000 ;
        RECT 4.265000 1.235000 4.455000 1.745000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.095000  0.085000  0.425000 1.040000 ;
      RECT 0.110000  1.825000  0.370000 2.905000 ;
      RECT 0.110000  2.905000  2.110000 3.075000 ;
      RECT 0.955000  0.085000  1.285000 0.685000 ;
      RECT 1.040000  1.960000  1.230000 2.905000 ;
      RECT 1.815000  0.085000  2.145000 0.645000 ;
      RECT 1.900000  2.105000  5.130000 2.285000 ;
      RECT 1.900000  2.285000  2.110000 2.905000 ;
      RECT 2.280000  2.455000  2.610000 3.245000 ;
      RECT 2.350000  0.255000  6.140000 0.425000 ;
      RECT 2.350000  0.425000  3.470000 0.645000 ;
      RECT 2.780000  2.285000  2.990000 3.075000 ;
      RECT 3.160000  2.465000  3.830000 3.245000 ;
      RECT 4.000000  2.285000  4.330000 3.075000 ;
      RECT 4.150000  0.425000  4.480000 0.895000 ;
      RECT 4.500000  2.455000  4.720000 3.245000 ;
      RECT 4.650000  0.595000  4.900000 0.815000 ;
      RECT 4.650000  0.815000  8.035000 0.985000 ;
      RECT 4.650000  0.985000  7.175000 1.025000 ;
      RECT 4.860000  1.755000 10.170000 1.925000 ;
      RECT 4.860000  1.925000  5.130000 2.105000 ;
      RECT 4.890000  2.285000  5.130000 3.075000 ;
      RECT 5.070000  0.425000  6.140000 0.645000 ;
      RECT 5.370000  2.105000  5.700000 3.245000 ;
      RECT 5.880000  1.925000  6.140000 3.075000 ;
      RECT 6.310000  2.105000  6.640000 3.245000 ;
      RECT 6.475000  0.255000  8.395000 0.425000 ;
      RECT 6.475000  0.425000  6.675000 0.645000 ;
      RECT 6.810000  1.925000  7.000000 3.075000 ;
      RECT 6.845000  0.615000  7.175000 0.815000 ;
      RECT 6.845000  1.025000  7.175000 1.145000 ;
      RECT 7.170000  2.105000  8.020000 3.245000 ;
      RECT 7.345000  0.425000  7.535000 0.645000 ;
      RECT 7.705000  0.615000  8.035000 0.815000 ;
      RECT 7.705000  0.985000  8.035000 1.145000 ;
      RECT 8.190000  1.925000  8.380000 3.075000 ;
      RECT 8.215000  0.425000  8.395000 0.860000 ;
      RECT 8.215000  0.860000 10.185000 1.030000 ;
      RECT 8.550000  2.105000  8.880000 3.245000 ;
      RECT 8.565000  0.085000  8.895000 0.690000 ;
      RECT 9.050000  1.925000  9.240000 3.075000 ;
      RECT 9.065000  0.315000  9.255000 0.860000 ;
      RECT 9.410000  2.105000  9.740000 3.245000 ;
      RECT 9.425000  0.085000  9.755000 0.690000 ;
      RECT 9.910000  1.925000 10.170000 3.075000 ;
      RECT 9.925000  0.315000 10.185000 0.860000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__a41oi_4
END LIBRARY
