* File: sky130_fd_sc_lp__o311ai_m.spice
* Created: Fri Aug 28 11:15:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o311ai_m  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_A_136_82#_M1008_d N_A1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_136_82#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_136_82#_M1004_d N_A3_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1006 A_394_82# N_B1_M1006_g N_A_136_82#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g A_394_82# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 A_148_403# N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1575 PD=0.63 PS=1.59 NRD=23.443 NRS=51.5943 M=1 R=2.8
+ SA=75000.3 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1001 A_220_403# N_A2_M1001_g A_148_403# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A3_M1002_g A_220_403# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.100375 AS=0.0588 PD=0.915 PS=0.7 NRD=39.8531 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.100375 PD=1.37 PS=0.915 NRD=0 NRS=39.8531 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.0799 P=10.25
c_38 VNB 0 3.15786e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o311ai_m.pxi.spice"
*
.ends
*
*
