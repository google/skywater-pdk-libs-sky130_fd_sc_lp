* File: sky130_fd_sc_lp__o2bb2ai_2.pex.spice
* Created: Fri Aug 28 11:12:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%A1_N 3 7 11 14 16 20 21 23 28 29 33
c84 21 0 1.2355e-19 $X=1.86 $Y=1.46
c85 14 0 1.36675e-19 $X=1.84 $Y=2.465
r86 28 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.51
+ $X2=0.46 $Y2=1.675
r87 28 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.46 $Y=1.51
+ $X2=0.46 $Y2=1.345
r88 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=1.51 $X2=0.46 $Y2=1.51
r89 23 40 5.64815 $w=7.18e-07 $l=3.4e-07 $layer=LI1_cond $X=0.445 $Y=1.665
+ $X2=0.445 $Y2=2.005
r90 23 29 2.57489 $w=7.18e-07 $l=1.55e-07 $layer=LI1_cond $X=0.445 $Y=1.665
+ $X2=0.445 $Y2=1.51
r91 21 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.46
+ $X2=1.86 $Y2=1.625
r92 21 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.46
+ $X2=1.86 $Y2=1.295
r93 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.86
+ $Y=1.46 $X2=1.86 $Y2=1.46
r94 18 20 16.8293 $w=3.13e-07 $l=4.6e-07 $layer=LI1_cond $X=1.852 $Y=1.92
+ $X2=1.852 $Y2=1.46
r95 17 40 9.50744 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=0.805 $Y=2.005
+ $X2=0.445 $Y2=2.005
r96 16 18 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=1.695 $Y=2.005
+ $X2=1.852 $Y2=1.92
r97 16 17 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=1.695 $Y=2.005
+ $X2=0.805 $Y2=2.005
r98 14 34 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.84 $Y=2.465
+ $X2=1.84 $Y2=1.625
r99 11 33 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.84 $Y=0.765
+ $X2=1.84 $Y2=1.295
r100 7 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.55 $Y=2.465
+ $X2=0.55 $Y2=1.675
r101 3 30 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.55 $Y=0.765
+ $X2=0.55 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%A2_N 1 3 6 8 10 13 15 16 24
c50 15 0 1.36675e-19 $X=1.2 $Y=1.295
r51 22 24 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.15 $Y=1.46
+ $X2=1.41 $Y2=1.46
r52 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.46 $X2=1.15 $Y2=1.46
r53 19 22 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.98 $Y=1.46
+ $X2=1.15 $Y2=1.46
r54 16 23 5.21694 $w=4.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.46
r55 15 23 4.199 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=1.295
+ $X2=1.22 $Y2=1.46
r56 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.625
+ $X2=1.41 $Y2=1.46
r57 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.41 $Y=1.625
+ $X2=1.41 $Y2=2.465
r58 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.46
r59 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=0.765
r60 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.625
+ $X2=0.98 $Y2=1.46
r61 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.98 $Y=1.625 $X2=0.98
+ $Y2=2.465
r62 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.295
+ $X2=0.98 $Y2=1.46
r63 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.98 $Y=1.295 $X2=0.98
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%A_125_367# 1 2 3 10 12 14 17 19 21 23 26
+ 28 29 32 34 40 42 45 47 49 51 55 58
c109 58 0 1.88051e-19 $X=2.4 $Y=1.37
c110 51 0 1.2355e-19 $X=1.625 $Y=2.345
r111 56 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.4 $Y=1.46 $X2=2.4
+ $Y2=1.37
r112 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=1.46 $X2=2.4 $Y2=1.46
r113 52 55 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=2.265 $Y=1.5
+ $X2=2.4 $Y2=1.5
r114 46 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=1.625
+ $X2=2.265 $Y2=1.5
r115 46 47 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.265 $Y=1.625
+ $X2=2.265 $Y2=2.26
r116 45 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=1.375
+ $X2=2.265 $Y2=1.5
r117 44 45 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.265 $Y=1.04
+ $X2=2.265 $Y2=1.375
r118 43 51 6.19399 $w=1.8e-07 $l=1.13e-07 $layer=LI1_cond $X=1.755 $Y=2.355
+ $X2=1.642 $Y2=2.355
r119 42 47 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.18 $Y=2.355
+ $X2=2.265 $Y2=2.26
r120 42 43 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=2.18 $Y=2.355
+ $X2=1.755 $Y2=2.355
r121 38 51 0.552779 $w=2.25e-07 $l=9.5e-08 $layer=LI1_cond $X=1.642 $Y=2.45
+ $X2=1.642 $Y2=2.355
r122 38 40 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=1.642 $Y=2.45
+ $X2=1.642 $Y2=2.91
r123 34 44 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.18 $Y=0.935
+ $X2=2.265 $Y2=1.04
r124 34 36 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=2.18 $Y=0.935
+ $X2=1.195 $Y2=0.935
r125 33 49 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.86 $Y=2.345
+ $X2=0.765 $Y2=2.345
r126 32 51 6.19399 $w=1.8e-07 $l=1.16893e-07 $layer=LI1_cond $X=1.53 $Y=2.345
+ $X2=1.642 $Y2=2.355
r127 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.53 $Y=2.345
+ $X2=0.86 $Y2=2.345
r128 24 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.28 $Y=1.445
+ $X2=3.28 $Y2=1.37
r129 24 26 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.28 $Y=1.445
+ $X2=3.28 $Y2=2.465
r130 21 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.28 $Y=1.295
+ $X2=3.28 $Y2=1.37
r131 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.28 $Y=1.295
+ $X2=3.28 $Y2=0.765
r132 20 28 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.925 $Y=1.37 $X2=2.85
+ $Y2=1.37
r133 19 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.205 $Y=1.37
+ $X2=3.28 $Y2=1.37
r134 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.205 $Y=1.37
+ $X2=2.925 $Y2=1.37
r135 15 28 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.85 $Y=1.445 $X2=2.85
+ $Y2=1.37
r136 15 17 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.85 $Y=1.445
+ $X2=2.85 $Y2=2.465
r137 12 28 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.85 $Y=1.295 $X2=2.85
+ $Y2=1.37
r138 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.85 $Y=1.295
+ $X2=2.85 $Y2=0.765
r139 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.565 $Y=1.37
+ $X2=2.4 $Y2=1.37
r140 10 28 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.775 $Y=1.37 $X2=2.85
+ $Y2=1.37
r141 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.775 $Y=1.37
+ $X2=2.565 $Y2=1.37
r142 3 51 600 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.345
r143 3 40 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.91
r144 2 49 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=0.625
+ $Y=1.835 $X2=0.765 $Y2=2.425
r145 1 36 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=1.055
+ $Y=0.345 $X2=1.195 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%B1 3 7 9 11 14 17 20 21 23 24 26 29 30
c84 30 0 1.48238e-19 $X=5.49 $Y=1.46
r85 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.46 $X2=5.49 $Y2=1.46
r86 26 30 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=5.5 $Y=1.665
+ $X2=5.5 $Y2=1.46
r87 25 26 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.5 $Y=1.92 $X2=5.5
+ $Y2=1.665
r88 23 25 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.325 $Y=2.005
+ $X2=5.5 $Y2=1.92
r89 23 24 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=5.325 $Y=2.005
+ $X2=3.815 $Y2=2.005
r90 21 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.51
+ $X2=3.73 $Y2=1.675
r91 21 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.51
+ $X2=3.73 $Y2=1.345
r92 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.51 $X2=3.73 $Y2=1.51
r93 18 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.69 $Y=1.92
+ $X2=3.815 $Y2=2.005
r94 18 20 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.69 $Y=1.92
+ $X2=3.69 $Y2=1.51
r95 16 29 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=5.155 $Y=1.46
+ $X2=5.49 $Y2=1.46
r96 16 17 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.155 $Y=1.46
+ $X2=5.08 $Y2=1.46
r97 12 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.08 $Y=1.625
+ $X2=5.08 $Y2=1.46
r98 12 14 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.08 $Y=1.625
+ $X2=5.08 $Y2=2.465
r99 9 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.08 $Y=1.295
+ $X2=5.08 $Y2=1.46
r100 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.08 $Y=1.295
+ $X2=5.08 $Y2=0.765
r101 7 33 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.79 $Y=0.765
+ $X2=3.79 $Y2=1.345
r102 3 34 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.75 $Y=2.465
+ $X2=3.75 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%B2 3 5 7 8 10 13 15 17 19 33
c56 33 0 1.48238e-19 $X=4.65 $Y=1.46
r57 31 33 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.61 $Y=1.46 $X2=4.65
+ $Y2=1.46
r58 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.61
+ $Y=1.46 $X2=4.61 $Y2=1.46
r59 29 31 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.22 $Y=1.46
+ $X2=4.61 $Y2=1.46
r60 27 29 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.18 $Y=1.46 $X2=4.22
+ $Y2=1.46
r61 19 32 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=5.04 $Y=1.48
+ $X2=4.61 $Y2=1.48
r62 17 32 1.10748 $w=5.38e-07 $l=5e-08 $layer=LI1_cond $X=4.56 $Y=1.48 $X2=4.61
+ $Y2=1.48
r63 15 17 10.6318 $w=5.38e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.48
+ $X2=4.56 $Y2=1.48
r64 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.65 $Y=1.625
+ $X2=4.65 $Y2=1.46
r65 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.65 $Y=1.625
+ $X2=4.65 $Y2=2.465
r66 8 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.65 $Y=1.295
+ $X2=4.65 $Y2=1.46
r67 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.65 $Y=1.295
+ $X2=4.65 $Y2=0.765
r68 5 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.22 $Y=1.295
+ $X2=4.22 $Y2=1.46
r69 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.22 $Y=1.295 $X2=4.22
+ $Y2=0.765
r70 1 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.18 $Y=1.625
+ $X2=4.18 $Y2=1.46
r71 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.18 $Y=1.625 $X2=4.18
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%VPWR 1 2 3 4 5 16 18 22 26 30 34 36 37 38
+ 39 41 51 62 67 71 78 80
r94 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r95 76 78 10.2749 $w=7.93e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=3.017 $X2=2.73
+ $Y2=3.017
r96 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 74 76 0.0752251 $w=7.93e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=3.017
+ $X2=2.64 $Y2=3.017
r98 70 71 10.8767 $w=7.93e-07 $l=1.3e-07 $layer=LI1_cond $X=2.055 $Y=3.017
+ $X2=1.925 $Y2=3.017
r99 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r100 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r102 59 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r103 59 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r105 56 80 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=3.515 $Y2=3.33
r106 56 58 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 55 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 54 78 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.73 $Y2=3.33
r109 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 51 80 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.4 $Y=3.33
+ $X2=3.515 $Y2=3.33
r111 51 54 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 50 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 50 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 49 71 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.925 $Y2=3.33
r115 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 47 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=3.33
+ $X2=1.195 $Y2=3.33
r117 47 49 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 45 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 45 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r120 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 42 64 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=3.33 $X2=0.25
+ $Y2=3.33
r122 42 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 41 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.195 $Y2=3.33
r124 41 44 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 39 55 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 39 77 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 37 58 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.13 $Y=3.33 $X2=5.04
+ $Y2=3.33
r128 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=3.33
+ $X2=5.295 $Y2=3.33
r129 36 61 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=5.46 $Y=3.33 $X2=5.52
+ $Y2=3.33
r130 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=3.33
+ $X2=5.295 $Y2=3.33
r131 32 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.295 $Y=3.245
+ $X2=5.295 $Y2=3.33
r132 32 34 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=5.295 $Y=3.245
+ $X2=5.295 $Y2=2.365
r133 28 80 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.245
+ $X2=3.515 $Y2=3.33
r134 28 30 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.515 $Y=3.245
+ $X2=3.515 $Y2=2.925
r135 24 74 0.15045 $w=7.93e-07 $l=1e-08 $layer=LI1_cond $X=2.625 $Y=3.017
+ $X2=2.635 $Y2=3.017
r136 24 70 8.57566 $w=7.93e-07 $l=5.7e-07 $layer=LI1_cond $X=2.625 $Y=3.017
+ $X2=2.055 $Y2=3.017
r137 24 26 33.8009 $w=2.08e-07 $l=6.4e-07 $layer=LI1_cond $X=2.625 $Y=2.62
+ $X2=2.625 $Y2=1.98
r138 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=3.33
r139 20 22 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=2.725
r140 16 64 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.25 $Y2=3.33
r141 16 18 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.335 $Y2=2.375
r142 5 34 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=5.155
+ $Y=1.835 $X2=5.295 $Y2=2.365
r143 4 30 600 $w=1.7e-07 $l=1.16726e-06 $layer=licon1_PDIFF $count=1 $X=3.355
+ $Y=1.835 $X2=3.515 $Y2=2.925
r144 3 74 600 $w=1.7e-07 $l=1.45101e-06 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.635 $Y2=2.97
r145 3 70 600 $w=1.7e-07 $l=1.0176e-06 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.785
r146 3 26 300 $w=1.7e-07 $l=7.89177e-07 $layer=licon1_PDIFF $count=2 $X=1.915
+ $Y=1.835 $X2=2.635 $Y2=1.98
r147 2 22 600 $w=1.7e-07 $l=9.57445e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.835 $X2=1.195 $Y2=2.725
r148 1 18 300 $w=1.7e-07 $l=5.9925e-07 $layer=licon1_PDIFF $count=2 $X=0.21
+ $Y=1.835 $X2=0.335 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%Y 1 2 3 12 14 15 16 17 18 19 28
c43 28 0 1.88051e-19 $X=3.065 $Y=0.68
r44 19 43 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.065 $Y=2.775
+ $X2=3.065 $Y2=2.91
r45 19 39 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.065 $Y=2.775
+ $X2=3.065 $Y2=2.59
r46 18 26 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=2.425
+ $X2=3.065 $Y2=2.26
r47 18 39 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=2.425
+ $X2=3.065 $Y2=2.59
r48 17 26 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.065 $Y=1.96
+ $X2=3.065 $Y2=2.26
r49 16 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.065 $Y=1.665
+ $X2=3.065 $Y2=1.96
r50 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.065 $Y=1.295
+ $X2=3.065 $Y2=1.665
r51 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.065 $Y=0.925
+ $X2=3.065 $Y2=1.295
r52 14 28 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.065 $Y=0.925
+ $X2=3.065 $Y2=0.68
r53 10 18 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=2.425
+ $X2=3.065 $Y2=2.425
r54 10 12 41.3832 $w=3.28e-07 $l=1.185e-06 $layer=LI1_cond $X=3.23 $Y=2.425
+ $X2=4.415 $Y2=2.425
r55 3 12 600 $w=1.7e-07 $l=6.65207e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.835 $X2=4.415 $Y2=2.425
r56 2 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=2.91
r57 2 17 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=1.96
r58 1 28 91 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=2 $X=2.925
+ $Y=0.345 $X2=3.065 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%A_765_367# 1 2 7 13
r16 11 13 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.835 $Y=2.76
+ $X2=4.835 $Y2=2.425
r17 7 11 7.03439 $w=3.15e-07 $l=2.06649e-07 $layer=LI1_cond $X=4.72 $Y=2.917
+ $X2=4.835 $Y2=2.76
r18 7 9 27.622 $w=3.13e-07 $l=7.55e-07 $layer=LI1_cond $X=4.72 $Y=2.917
+ $X2=3.965 $Y2=2.917
r19 2 13 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=4.725
+ $Y=1.835 $X2=4.865 $Y2=2.425
r20 1 9 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=1.835 $X2=3.965 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%VGND 1 2 3 4 13 15 19 23 27 30 31 32 34 42
+ 52 53 59 62
r73 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r74 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r75 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r76 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r77 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r78 50 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r79 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r80 47 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.005
+ $Y2=0
r81 47 49 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.56
+ $Y2=0
r82 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r83 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r84 43 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.055
+ $Y2=0
r85 43 45 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.22 $Y=0 $X2=3.6
+ $Y2=0
r86 42 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=4.005
+ $Y2=0
r87 42 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r88 41 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r89 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r90 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r91 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r92 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r93 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r94 35 56 4.40897 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=0 $X2=0.237
+ $Y2=0
r95 35 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.475 $Y=0 $X2=0.72
+ $Y2=0
r96 34 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.055
+ $Y2=0
r97 34 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r98 32 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r99 32 60 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r100 30 49 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.7 $Y=0 $X2=4.56
+ $Y2=0
r101 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.7 $Y=0 $X2=4.865
+ $Y2=0
r102 29 52 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.03 $Y=0 $X2=5.52
+ $Y2=0
r103 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.03 $Y=0 $X2=4.865
+ $Y2=0
r104 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=0.085
+ $X2=4.865 $Y2=0
r105 25 27 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.865 $Y=0.085
+ $X2=4.865 $Y2=0.575
r106 21 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.005 $Y=0.085
+ $X2=4.005 $Y2=0
r107 21 23 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.005 $Y=0.085
+ $X2=4.005 $Y2=0.575
r108 17 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r109 17 19 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.535
r110 13 56 3.14927 $w=3.05e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.322 $Y=0.085
+ $X2=0.237 $Y2=0
r111 13 15 15.3029 $w=3.03e-07 $l=4.05e-07 $layer=LI1_cond $X=0.322 $Y=0.085
+ $X2=0.322 $Y2=0.49
r112 4 27 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=4.725
+ $Y=0.345 $X2=4.865 $Y2=0.575
r113 3 23 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=3.865
+ $Y=0.345 $X2=4.005 $Y2=0.575
r114 2 19 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.345 $X2=2.055 $Y2=0.535
r115 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.345 $X2=0.335 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%A_125_69# 1 2 7 9 13
r17 11 16 2.78134 $w=3.55e-07 $l=1.08e-07 $layer=LI1_cond $X=0.86 $Y=0.482
+ $X2=0.752 $Y2=0.482
r18 11 13 24.8343 $w=3.53e-07 $l=7.65e-07 $layer=LI1_cond $X=0.86 $Y=0.482
+ $X2=1.625 $Y2=0.482
r19 7 16 4.58406 $w=2.15e-07 $l=1.78e-07 $layer=LI1_cond $X=0.752 $Y=0.66
+ $X2=0.752 $Y2=0.482
r20 7 9 14.2045 $w=2.13e-07 $l=2.65e-07 $layer=LI1_cond $X=0.752 $Y=0.66
+ $X2=0.752 $Y2=0.925
r21 2 13 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.345 $X2=1.625 $Y2=0.495
r22 1 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.345 $X2=0.765 $Y2=0.47
r23 1 9 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.345 $X2=0.765 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_2%A_502_69# 1 2 3 4 15 17 18 23 24 27 29 33
+ 36
r54 31 33 16.8434 $w=2.58e-07 $l=3.8e-07 $layer=LI1_cond $X=5.33 $Y=0.87
+ $X2=5.33 $Y2=0.49
r55 30 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.53 $Y=0.955
+ $X2=4.435 $Y2=0.955
r56 29 31 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.2 $Y=0.955
+ $X2=5.33 $Y2=0.87
r57 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.2 $Y=0.955
+ $X2=4.53 $Y2=0.955
r58 25 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.87
+ $X2=4.435 $Y2=0.955
r59 25 27 22.1818 $w=1.88e-07 $l=3.8e-07 $layer=LI1_cond $X=4.435 $Y=0.87
+ $X2=4.435 $Y2=0.49
r60 23 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.34 $Y=0.955
+ $X2=4.435 $Y2=0.955
r61 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.34 $Y=0.955
+ $X2=3.67 $Y2=0.955
r62 20 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.54 $Y=0.87
+ $X2=3.67 $Y2=0.955
r63 20 22 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=3.54 $Y=0.87 $X2=3.54
+ $Y2=0.47
r64 19 22 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=3.54 $Y=0.425
+ $X2=3.54 $Y2=0.47
r65 17 19 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.41 $Y=0.34
+ $X2=3.54 $Y2=0.425
r66 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.41 $Y=0.34
+ $X2=2.73 $Y2=0.34
r67 13 18 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.625 $Y=0.425
+ $X2=2.73 $Y2=0.34
r68 13 15 3.4329 $w=2.08e-07 $l=6.5e-08 $layer=LI1_cond $X=2.625 $Y=0.425
+ $X2=2.625 $Y2=0.49
r69 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.155
+ $Y=0.345 $X2=5.295 $Y2=0.49
r70 3 36 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=4.295
+ $Y=0.345 $X2=4.435 $Y2=0.955
r71 3 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.295
+ $Y=0.345 $X2=4.435 $Y2=0.49
r72 2 22 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=3.355
+ $Y=0.345 $X2=3.535 $Y2=0.47
r73 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.51
+ $Y=0.345 $X2=2.635 $Y2=0.49
.ends

