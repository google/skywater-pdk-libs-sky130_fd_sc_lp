* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_800_473# a_809_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_587_47# a_371_473# a_659_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_41_464# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_371_473# a_249_70# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_659_47# a_249_70# a_767_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_809_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_809_21# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_371_473# a_249_70# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND GATE a_249_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_809_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_41_464# a_587_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR GATE a_249_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_809_21# a_659_47# a_1056_73# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_1056_73# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_659_47# a_371_473# a_800_473# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_767_47# a_809_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR a_659_47# a_809_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR a_41_464# a_623_473# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_623_473# a_249_70# a_659_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_41_464# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
