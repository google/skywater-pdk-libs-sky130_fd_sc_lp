* File: sky130_fd_sc_lp__mux2i_2.spice
* Created: Fri Aug 28 10:45:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2i_2.pex.spice"
.subckt sky130_fd_sc_lp__mux2i_2  VNB VPB S A0 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_S_M1012_g N_A_44_367#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1012_d N_A_44_367#_M1009_g N_A_251_47#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_A_44_367#_M1017_g N_A_251_47#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1017_d N_S_M1003_g N_A_423_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_S_M1010_g N_A_423_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_A0_M1001_g N_A_251_47#_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1013 N_Y_M1013_d N_A0_M1013_g N_A_251_47#_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_423_47#_M1007_d N_A1_M1007_g N_Y_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=11.424 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_A_423_47#_M1007_d N_A1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.2226 PD=1.2 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.7 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_S_M1006_g N_A_44_367#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2961 AS=0.3339 PD=1.73 PS=3.05 NRD=15.6221 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 N_A_251_367#_M1002_d N_A_44_367#_M1002_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.2961 PD=1.54 PS=1.73 NRD=0 NRS=14.0658 M=1 R=8.4
+ SA=75000.8 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1015 N_A_251_367#_M1002_d N_A_44_367#_M1015_g N_VPWR_M1015_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.290975 PD=1.54 PS=1.795 NRD=0 NRS=13.2778 M=1
+ R=8.4 SA=75001.2 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1004 N_A_455_367#_M1004_d N_S_M1004_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.290975 PD=1.54 PS=1.795 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75001.8
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1014 N_A_455_367#_M1004_d N_S_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.53155 PD=1.54 PS=3.51 NRD=0 NRS=18.7544 M=1 R=8.4 SA=75002.3
+ SB=75000.3 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A0_M1005_g N_A_455_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1011_d N_A0_M1011_g N_A_455_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1011_d N_A1_M1000_g N_A_251_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_Y_M1016_d N_A1_M1016_g N_A_251_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__mux2i_2.pxi.spice"
*
.ends
*
*
