* File: sky130_fd_sc_lp__o2111a_4.pxi.spice
* Created: Fri Aug 28 11:00:13 2020
* 
x_PM_SKY130_FD_SC_LP__O2111A_4%D1 N_D1_M1013_g N_D1_c_147_n N_D1_M1018_g
+ N_D1_M1026_g N_D1_c_149_n N_D1_M1021_g D1 N_D1_c_151_n
+ PM_SKY130_FD_SC_LP__O2111A_4%D1
x_PM_SKY130_FD_SC_LP__O2111A_4%C1 N_C1_M1016_g N_C1_M1007_g N_C1_M1027_g
+ N_C1_M1022_g N_C1_c_197_n N_C1_c_190_n N_C1_c_191_n N_C1_c_244_p N_C1_c_192_n
+ N_C1_c_193_n C1 PM_SKY130_FD_SC_LP__O2111A_4%C1
x_PM_SKY130_FD_SC_LP__O2111A_4%B1 N_B1_M1005_g N_B1_M1004_g N_B1_M1015_g
+ N_B1_M1017_g B1 N_B1_c_287_n N_B1_c_288_n PM_SKY130_FD_SC_LP__O2111A_4%B1
x_PM_SKY130_FD_SC_LP__O2111A_4%A2 N_A2_M1006_g N_A2_c_337_n N_A2_c_338_n
+ N_A2_M1019_g N_A2_c_349_n N_A2_M1024_g N_A2_c_339_n N_A2_c_340_n N_A2_M1023_g
+ N_A2_c_342_n N_A2_c_343_n N_A2_c_344_n A2 A2 N_A2_c_345_n N_A2_c_346_n A2
+ PM_SKY130_FD_SC_LP__O2111A_4%A2
x_PM_SKY130_FD_SC_LP__O2111A_4%A1 N_A1_c_462_n N_A1_M1001_g N_A1_c_453_n
+ N_A1_c_454_n N_A1_c_455_n N_A1_M1000_g N_A1_c_465_n N_A1_M1011_g N_A1_c_456_n
+ N_A1_c_457_n N_A1_M1008_g N_A1_c_458_n N_A1_c_459_n A1 A1 N_A1_c_461_n
+ PM_SKY130_FD_SC_LP__O2111A_4%A1
x_PM_SKY130_FD_SC_LP__O2111A_4%A_32_367# N_A_32_367#_M1018_s N_A_32_367#_M1013_s
+ N_A_32_367#_M1026_s N_A_32_367#_M1004_s N_A_32_367#_M1022_s
+ N_A_32_367#_M1024_s N_A_32_367#_M1003_g N_A_32_367#_M1002_g
+ N_A_32_367#_M1010_g N_A_32_367#_M1009_g N_A_32_367#_M1012_g
+ N_A_32_367#_M1014_g N_A_32_367#_M1020_g N_A_32_367#_M1025_g
+ N_A_32_367#_c_532_n N_A_32_367#_c_533_n N_A_32_367#_c_534_n
+ N_A_32_367#_c_535_n N_A_32_367#_c_629_p N_A_32_367#_c_562_n
+ N_A_32_367#_c_630_p N_A_32_367#_c_567_n N_A_32_367#_c_581_n
+ N_A_32_367#_c_536_n N_A_32_367#_c_537_n N_A_32_367#_c_525_n
+ N_A_32_367#_c_526_n N_A_32_367#_c_658_p N_A_32_367#_c_539_n
+ N_A_32_367#_c_572_n N_A_32_367#_c_573_n N_A_32_367#_c_540_n
+ N_A_32_367#_c_527_n PM_SKY130_FD_SC_LP__O2111A_4%A_32_367#
x_PM_SKY130_FD_SC_LP__O2111A_4%VPWR N_VPWR_M1013_d N_VPWR_M1016_d N_VPWR_M1017_d
+ N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_M1025_d N_VPWR_c_704_n
+ N_VPWR_c_705_n N_VPWR_c_706_n N_VPWR_c_707_n N_VPWR_c_708_n N_VPWR_c_709_n
+ N_VPWR_c_710_n N_VPWR_c_711_n N_VPWR_c_712_n N_VPWR_c_713_n VPWR
+ N_VPWR_c_714_n N_VPWR_c_715_n N_VPWR_c_716_n N_VPWR_c_717_n N_VPWR_c_718_n
+ N_VPWR_c_719_n N_VPWR_c_720_n N_VPWR_c_721_n N_VPWR_c_722_n N_VPWR_c_723_n
+ N_VPWR_c_724_n N_VPWR_c_703_n PM_SKY130_FD_SC_LP__O2111A_4%VPWR
x_PM_SKY130_FD_SC_LP__O2111A_4%A_741_367# N_A_741_367#_M1006_d
+ N_A_741_367#_M1011_d N_A_741_367#_c_824_n N_A_741_367#_c_829_n
+ N_A_741_367#_c_830_n PM_SKY130_FD_SC_LP__O2111A_4%A_741_367#
x_PM_SKY130_FD_SC_LP__O2111A_4%X N_X_M1003_s N_X_M1012_s N_X_M1002_s N_X_M1014_s
+ N_X_c_893_p N_X_c_879_n N_X_c_839_n N_X_c_840_n N_X_c_845_n N_X_c_846_n
+ N_X_c_894_p N_X_c_883_n N_X_c_841_n N_X_c_842_n N_X_c_847_n X X N_X_c_843_n X
+ PM_SKY130_FD_SC_LP__O2111A_4%X
x_PM_SKY130_FD_SC_LP__O2111A_4%A_32_65# N_A_32_65#_M1018_d N_A_32_65#_M1021_d
+ N_A_32_65#_M1027_s N_A_32_65#_c_899_n N_A_32_65#_c_900_n N_A_32_65#_c_901_n
+ N_A_32_65#_c_902_n N_A_32_65#_c_903_n N_A_32_65#_c_904_n
+ PM_SKY130_FD_SC_LP__O2111A_4%A_32_65#
x_PM_SKY130_FD_SC_LP__O2111A_4%A_289_65# N_A_289_65#_M1007_d N_A_289_65#_M1015_s
+ N_A_289_65#_c_948_n N_A_289_65#_c_950_n N_A_289_65#_c_951_n
+ N_A_289_65#_c_953_n PM_SKY130_FD_SC_LP__O2111A_4%A_289_65#
x_PM_SKY130_FD_SC_LP__O2111A_4%A_389_65# N_A_389_65#_M1005_d N_A_389_65#_M1019_d
+ N_A_389_65#_M1008_s N_A_389_65#_c_970_n N_A_389_65#_c_971_n
+ N_A_389_65#_c_972_n N_A_389_65#_c_973_n N_A_389_65#_c_1018_p
+ N_A_389_65#_c_989_n N_A_389_65#_c_990_n N_A_389_65#_c_994_n
+ N_A_389_65#_c_974_n N_A_389_65#_c_995_n PM_SKY130_FD_SC_LP__O2111A_4%A_389_65#
x_PM_SKY130_FD_SC_LP__O2111A_4%VGND N_VGND_M1019_s N_VGND_M1000_d N_VGND_M1023_s
+ N_VGND_M1010_d N_VGND_M1020_d N_VGND_c_1034_n N_VGND_c_1035_n N_VGND_c_1036_n
+ N_VGND_c_1037_n N_VGND_c_1038_n N_VGND_c_1039_n N_VGND_c_1040_n
+ N_VGND_c_1041_n N_VGND_c_1042_n VGND N_VGND_c_1043_n N_VGND_c_1044_n
+ N_VGND_c_1045_n N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n
+ N_VGND_c_1049_n PM_SKY130_FD_SC_LP__O2111A_4%VGND
cc_1 VNB N_D1_M1013_g 0.00373837f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_2 VNB N_D1_c_147_n 0.0197233f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.275
cc_3 VNB N_D1_M1026_g 0.00223111f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.465
cc_4 VNB N_D1_c_149_n 0.0159594f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.275
cc_5 VNB D1 0.0230591f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_D1_c_151_n 0.0711297f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.44
cc_7 VNB N_C1_M1007_g 0.0207719f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.745
cc_8 VNB N_C1_M1027_g 0.0236687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C1_c_190_n 0.0230662f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.44
cc_10 VNB N_C1_c_191_n 0.00359708f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.44
cc_11 VNB N_C1_c_192_n 0.00224737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C1_c_193_n 0.0325167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB C1 6.51408e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_M1005_g 0.0203934f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_15 VNB N_B1_M1015_g 0.0192059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_287_n 0.00165125f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.44
cc_17 VNB N_B1_c_288_n 0.0316108f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_18 VNB N_A2_M1006_g 0.00732257f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_19 VNB N_A2_c_337_n 0.0200807f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.275
cc_20 VNB N_A2_c_338_n 0.0196339f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.745
cc_21 VNB N_A2_c_339_n 0.00550934f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.745
cc_22 VNB N_A2_c_340_n 0.00580369f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.745
cc_23 VNB N_A2_M1023_g 0.0233915f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.44
cc_24 VNB N_A2_c_342_n 0.0120426f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.44
cc_25 VNB N_A2_c_343_n 0.00811388f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.44
cc_26 VNB N_A2_c_344_n 0.025636f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_27 VNB N_A2_c_345_n 0.0374704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_c_346_n 0.00421826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB A2 0.00540502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_453_n 0.00622884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A1_c_454_n 0.00475252f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.275
cc_32 VNB N_A1_c_455_n 0.0151292f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.745
cc_33 VNB N_A1_c_456_n 0.017468f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.275
cc_34 VNB N_A1_c_457_n 0.0151292f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.745
cc_35 VNB N_A1_c_458_n 0.00995517f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.44
cc_36 VNB N_A1_c_459_n 0.00361415f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.44
cc_37 VNB A1 0.00749364f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.44
cc_38 VNB N_A1_c_461_n 0.0194502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_32_367#_M1003_g 0.0242861f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.44
cc_40 VNB N_A_32_367#_M1010_g 0.0217542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_32_367#_M1012_g 0.0217337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_32_367#_M1020_g 0.0265001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_32_367#_c_525_n 6.66824e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_32_367#_c_526_n 0.00183575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_32_367#_c_527_n 0.0782818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VPWR_c_703_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_X_c_839_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.44
cc_48 VNB N_X_c_840_n 0.00368316f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_49 VNB N_X_c_841_n 0.00108129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_X_c_842_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_X_c_843_n 0.0142938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB X 0.0190659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_32_65#_c_899_n 0.023066f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.275
cc_54 VNB N_A_32_65#_c_900_n 0.00464669f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.745
cc_55 VNB N_A_32_65#_c_901_n 0.00925098f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_56 VNB N_A_32_65#_c_902_n 0.0225009f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.44
cc_57 VNB N_A_32_65#_c_903_n 0.00342074f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.44
cc_58 VNB N_A_32_65#_c_904_n 0.00953706f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_59 VNB N_A_289_65#_c_948_n 0.00272872f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.465
cc_60 VNB N_A_389_65#_c_970_n 0.0168771f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.465
cc_61 VNB N_A_389_65#_c_971_n 0.00761485f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.745
cc_62 VNB N_A_389_65#_c_972_n 0.00432904f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.745
cc_63 VNB N_A_389_65#_c_973_n 0.00447686f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_64 VNB N_A_389_65#_c_974_n 0.00200998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1034_n 0.00450232f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.44
cc_66 VNB N_VGND_c_1035_n 0.0135029f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.44
cc_67 VNB N_VGND_c_1036_n 3.27005e-19 $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_68 VNB N_VGND_c_1037_n 0.00395069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1038_n 3.15212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1039_n 0.0146719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1040_n 0.0277511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1041_n 0.0891592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1042_n 0.00468472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1043_n 0.0148035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1044_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1045_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1046_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1047_n 0.00509388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1048_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1049_n 0.396253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VPB N_D1_M1013_g 0.0264218f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_82 VPB N_D1_M1026_g 0.0189989f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.465
cc_83 VPB N_C1_M1016_g 0.0192726f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_84 VPB N_C1_M1022_g 0.0239397f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_85 VPB N_C1_c_197_n 0.00129713f $X=-0.19 $Y=1.655 $X2=0.285 $Y2=1.44
cc_86 VPB N_C1_c_190_n 0.0064305f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=1.44
cc_87 VPB N_C1_c_193_n 0.00945627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB C1 0.0013035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_B1_M1004_g 0.0188619f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.745
cc_90 VPB N_B1_M1017_g 0.0183525f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_91 VPB N_B1_c_287_n 0.00365255f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.44
cc_92 VPB N_B1_c_288_n 0.00471481f $X=-0.19 $Y=1.655 $X2=0.237 $Y2=1.295
cc_93 VPB N_A2_M1006_g 0.0256679f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_94 VPB N_A2_c_349_n 0.0203257f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.465
cc_95 VPB N_A2_c_339_n 0.0048066f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=0.745
cc_96 VPB N_A2_c_340_n 0.00229348f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=0.745
cc_97 VPB N_A2_c_344_n 0.0118685f $X=-0.19 $Y=1.655 $X2=0.237 $Y2=1.295
cc_98 VPB A2 0.004158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A1_c_462_n 0.0159151f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.605
cc_100 VPB N_A1_c_453_n 0.00351058f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A1_c_454_n 0.00204574f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=1.275
cc_102 VPB N_A1_c_465_n 0.0159089f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.465
cc_103 VPB N_A1_c_459_n 0.00573162f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.44
cc_104 VPB A1 0.00680951f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.44
cc_105 VPB N_A_32_367#_M1002_g 0.0224981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_32_367#_M1009_g 0.0188385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_32_367#_M1014_g 0.0188385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_32_367#_M1025_g 0.0231294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_32_367#_c_532_n 0.00897476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_32_367#_c_533_n 0.0412714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_32_367#_c_534_n 4.07949e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_32_367#_c_535_n 7.99442e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_32_367#_c_536_n 0.00933283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_32_367#_c_537_n 0.0168272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_32_367#_c_525_n 0.00110952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_32_367#_c_539_n 0.00519241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_32_367#_c_540_n 0.00585173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_32_367#_c_527_n 0.010874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_704_n 4.05231e-19 $X=-0.19 $Y=1.655 $X2=0.237 $Y2=1.295
cc_120 VPB N_VPWR_c_705_n 0.00432043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_706_n 4.06898e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_707_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_708_n 0.0124894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_709_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_710_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_711_n 0.0415892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_712_n 0.034712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_713_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_714_n 0.0161714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_715_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_716_n 0.0149824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_717_n 0.0282439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_718_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_719_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_720_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_721_n 0.00628274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_722_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_723_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_724_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_703_n 0.0563694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_X_c_845_n 0.00304705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_X_c_846_n 0.00202714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_X_c_847_n 0.011898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB X 0.00528999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 N_D1_M1026_g N_C1_M1016_g 0.0182301f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_146 N_D1_c_149_n N_C1_M1007_g 0.0202361f $X=0.94 $Y=1.275 $X2=0 $Y2=0
cc_147 N_D1_M1026_g N_C1_c_197_n 5.22957e-19 $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_148 N_D1_c_151_n N_C1_c_190_n 0.0209203f $X=0.93 $Y=1.44 $X2=0 $Y2=0
cc_149 N_D1_c_151_n N_C1_c_191_n 9.19637e-19 $X=0.93 $Y=1.44 $X2=0 $Y2=0
cc_150 D1 N_A_32_367#_c_532_n 0.0190206f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_151 N_D1_c_151_n N_A_32_367#_c_532_n 0.00200427f $X=0.93 $Y=1.44 $X2=0 $Y2=0
cc_152 N_D1_M1013_g N_A_32_367#_c_534_n 0.0140124f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_153 D1 N_A_32_367#_c_534_n 5.54955e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_154 N_D1_c_151_n N_A_32_367#_c_534_n 0.00135357f $X=0.93 $Y=1.44 $X2=0 $Y2=0
cc_155 N_D1_M1013_g N_A_32_367#_c_535_n 0.0114484f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_156 N_D1_c_147_n N_A_32_367#_c_535_n 0.0144186f $X=0.51 $Y=1.275 $X2=0 $Y2=0
cc_157 N_D1_M1026_g N_A_32_367#_c_535_n 0.00626716f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_158 N_D1_c_149_n N_A_32_367#_c_535_n 0.00862508f $X=0.94 $Y=1.275 $X2=0 $Y2=0
cc_159 D1 N_A_32_367#_c_535_n 0.02969f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_160 N_D1_c_151_n N_A_32_367#_c_535_n 0.0234132f $X=0.93 $Y=1.44 $X2=0 $Y2=0
cc_161 N_D1_M1013_g N_A_32_367#_c_539_n 0.00243252f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_162 N_D1_M1026_g N_A_32_367#_c_539_n 0.0156297f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_163 N_D1_c_151_n N_A_32_367#_c_539_n 7.31956e-19 $X=0.93 $Y=1.44 $X2=0 $Y2=0
cc_164 N_D1_M1013_g N_VPWR_c_704_n 0.01556f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_165 N_D1_M1026_g N_VPWR_c_704_n 0.0136735f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_166 N_D1_M1013_g N_VPWR_c_714_n 0.00486043f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_167 N_D1_M1026_g N_VPWR_c_715_n 0.00486043f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_168 N_D1_M1013_g N_VPWR_c_703_n 0.00920269f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_169 N_D1_M1026_g N_VPWR_c_703_n 0.0082726f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_170 D1 N_A_32_65#_c_899_n 0.0223247f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_171 N_D1_c_151_n N_A_32_65#_c_899_n 0.00169228f $X=0.93 $Y=1.44 $X2=0 $Y2=0
cc_172 N_D1_c_147_n N_A_32_65#_c_900_n 0.0125027f $X=0.51 $Y=1.275 $X2=0 $Y2=0
cc_173 N_D1_c_149_n N_A_32_65#_c_900_n 0.0118056f $X=0.94 $Y=1.275 $X2=0 $Y2=0
cc_174 N_D1_c_149_n N_A_32_65#_c_903_n 7.38449e-19 $X=0.94 $Y=1.275 $X2=0 $Y2=0
cc_175 N_D1_c_147_n N_VGND_c_1041_n 0.00302501f $X=0.51 $Y=1.275 $X2=0 $Y2=0
cc_176 N_D1_c_149_n N_VGND_c_1041_n 0.00302501f $X=0.94 $Y=1.275 $X2=0 $Y2=0
cc_177 N_D1_c_147_n N_VGND_c_1049_n 0.00471752f $X=0.51 $Y=1.275 $X2=0 $Y2=0
cc_178 N_D1_c_149_n N_VGND_c_1049_n 0.00435646f $X=0.94 $Y=1.275 $X2=0 $Y2=0
cc_179 N_C1_M1007_g N_B1_M1005_g 0.0269332f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_180 N_C1_M1016_g N_B1_M1004_g 0.0368493f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_181 N_C1_c_197_n N_B1_M1004_g 0.00352765f $X=1.515 $Y=1.95 $X2=0 $Y2=0
cc_182 C1 N_B1_M1004_g 0.0108535f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_183 N_C1_M1027_g N_B1_M1015_g 0.0341794f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_184 N_C1_M1022_g N_B1_M1017_g 0.0341794f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_185 C1 N_B1_M1017_g 0.0104125f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_186 N_C1_M1016_g N_B1_c_287_n 2.96755e-19 $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_187 N_C1_c_197_n N_B1_c_287_n 0.0112396f $X=1.515 $Y=1.95 $X2=0 $Y2=0
cc_188 N_C1_c_190_n N_B1_c_287_n 8.36565e-19 $X=1.39 $Y=1.51 $X2=0 $Y2=0
cc_189 N_C1_c_191_n N_B1_c_287_n 0.0192814f $X=1.515 $Y=1.535 $X2=0 $Y2=0
cc_190 N_C1_c_192_n N_B1_c_287_n 0.0136574f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_191 N_C1_c_193_n N_B1_c_287_n 3.75387e-19 $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_192 C1 N_B1_c_287_n 0.054488f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_193 N_C1_c_197_n N_B1_c_288_n 4.19116e-19 $X=1.515 $Y=1.95 $X2=0 $Y2=0
cc_194 N_C1_c_190_n N_B1_c_288_n 0.0193006f $X=1.39 $Y=1.51 $X2=0 $Y2=0
cc_195 N_C1_c_191_n N_B1_c_288_n 7.07677e-19 $X=1.515 $Y=1.535 $X2=0 $Y2=0
cc_196 N_C1_c_192_n N_B1_c_288_n 0.00122101f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_197 N_C1_c_193_n N_B1_c_288_n 0.0341794f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_198 C1 N_B1_c_288_n 0.00515467f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_199 N_C1_c_193_n N_A2_M1006_g 0.00331913f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_200 N_C1_M1027_g N_A2_c_345_n 0.00197109f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_201 N_C1_c_193_n N_A2_c_345_n 0.0053224f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_202 N_C1_M1027_g N_A2_c_346_n 5.34529e-19 $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_203 N_C1_M1027_g A2 0.00158813f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_204 N_C1_M1022_g A2 0.00114774f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_205 N_C1_c_192_n A2 0.00751168f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_206 N_C1_c_193_n A2 0.00439253f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_207 C1 A2 0.00440378f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_208 C1 N_A_32_367#_M1004_s 0.00333507f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_209 N_C1_M1016_g N_A_32_367#_c_535_n 4.20018e-19 $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_210 N_C1_M1007_g N_A_32_367#_c_535_n 5.2411e-19 $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_211 N_C1_c_197_n N_A_32_367#_c_535_n 0.00469119f $X=1.515 $Y=1.95 $X2=0 $Y2=0
cc_212 N_C1_c_190_n N_A_32_367#_c_535_n 7.82328e-19 $X=1.39 $Y=1.51 $X2=0 $Y2=0
cc_213 N_C1_c_191_n N_A_32_367#_c_535_n 0.0095987f $X=1.515 $Y=1.535 $X2=0 $Y2=0
cc_214 N_C1_M1016_g N_A_32_367#_c_562_n 0.0152376f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_215 N_C1_c_190_n N_A_32_367#_c_562_n 2.87136e-19 $X=1.39 $Y=1.51 $X2=0 $Y2=0
cc_216 N_C1_c_191_n N_A_32_367#_c_562_n 0.00343528f $X=1.515 $Y=1.535 $X2=0
+ $Y2=0
cc_217 N_C1_c_244_p N_A_32_367#_c_562_n 0.00882278f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_218 C1 N_A_32_367#_c_562_n 0.0201202f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_219 N_C1_M1022_g N_A_32_367#_c_567_n 0.0123944f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_220 C1 N_A_32_367#_c_567_n 0.0283894f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_221 N_C1_c_197_n N_A_32_367#_c_539_n 0.00513045f $X=1.515 $Y=1.95 $X2=0 $Y2=0
cc_222 N_C1_c_190_n N_A_32_367#_c_539_n 5.80622e-19 $X=1.39 $Y=1.51 $X2=0 $Y2=0
cc_223 N_C1_c_191_n N_A_32_367#_c_539_n 0.0018223f $X=1.515 $Y=1.535 $X2=0 $Y2=0
cc_224 C1 N_A_32_367#_c_572_n 0.0135055f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_225 N_C1_c_192_n N_A_32_367#_c_573_n 0.00375366f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_226 N_C1_c_193_n N_A_32_367#_c_573_n 0.00578893f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_227 C1 N_A_32_367#_c_573_n 0.0164008f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_228 N_C1_c_197_n N_VPWR_M1016_d 0.00134539f $X=1.515 $Y=1.95 $X2=0 $Y2=0
cc_229 N_C1_c_244_p N_VPWR_M1016_d 0.00117408f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_230 C1 N_VPWR_M1016_d 0.0066872f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_231 C1 N_VPWR_M1017_d 0.00775772f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_232 N_C1_M1016_g N_VPWR_c_704_n 6.3841e-19 $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_233 N_C1_M1016_g N_VPWR_c_705_n 0.00262861f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_234 N_C1_M1022_g N_VPWR_c_706_n 0.0118283f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_235 N_C1_M1022_g N_VPWR_c_712_n 0.00486043f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_236 N_C1_M1016_g N_VPWR_c_715_n 0.00585385f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_237 N_C1_M1016_g N_VPWR_c_703_n 0.0108771f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_238 N_C1_M1022_g N_VPWR_c_703_n 0.00588233f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_239 N_C1_M1007_g N_A_32_65#_c_900_n 8.31364e-19 $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_240 N_C1_M1007_g N_A_32_65#_c_902_n 0.0133991f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_241 N_C1_M1027_g N_A_32_65#_c_902_n 0.0136051f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_242 N_C1_c_190_n N_A_32_65#_c_902_n 0.00386072f $X=1.39 $Y=1.51 $X2=0 $Y2=0
cc_243 N_C1_c_191_n N_A_32_65#_c_902_n 0.0250888f $X=1.515 $Y=1.535 $X2=0 $Y2=0
cc_244 N_C1_c_192_n N_A_32_65#_c_902_n 0.0317408f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_245 N_C1_c_193_n N_A_32_65#_c_902_n 0.00773881f $X=2.82 $Y=1.51 $X2=0 $Y2=0
cc_246 N_C1_c_190_n N_A_32_65#_c_903_n 6.41898e-19 $X=1.39 $Y=1.51 $X2=0 $Y2=0
cc_247 N_C1_c_191_n N_A_32_65#_c_903_n 0.00205129f $X=1.515 $Y=1.535 $X2=0 $Y2=0
cc_248 N_C1_M1007_g N_A_289_65#_c_948_n 0.00508387f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_249 N_C1_M1007_g N_A_289_65#_c_950_n 0.00226088f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_250 N_C1_M1027_g N_A_289_65#_c_951_n 0.0032337f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_251 N_C1_M1027_g N_A_389_65#_c_970_n 0.0132977f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_252 N_C1_M1027_g N_A_389_65#_c_971_n 0.00406574f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_253 N_C1_M1027_g N_A_389_65#_c_974_n 7.15369e-19 $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_254 N_C1_M1007_g N_VGND_c_1041_n 0.0046877f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_255 N_C1_M1027_g N_VGND_c_1041_n 0.00302501f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_256 N_C1_M1007_g N_VGND_c_1049_n 0.00909832f $X=1.37 $Y=0.745 $X2=0 $Y2=0
cc_257 N_C1_M1027_g N_VGND_c_1049_n 0.00485634f $X=2.73 $Y=0.745 $X2=0 $Y2=0
cc_258 N_B1_M1004_g N_A_32_367#_c_562_n 0.0133747f $X=1.87 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B1_M1017_g N_A_32_367#_c_567_n 0.00999655f $X=2.3 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B1_M1004_g N_VPWR_c_705_n 0.0025782f $X=1.87 $Y=2.465 $X2=0 $Y2=0
cc_261 N_B1_M1004_g N_VPWR_c_706_n 5.9121e-19 $X=1.87 $Y=2.465 $X2=0 $Y2=0
cc_262 N_B1_M1017_g N_VPWR_c_706_n 0.0102609f $X=2.3 $Y=2.465 $X2=0 $Y2=0
cc_263 N_B1_M1004_g N_VPWR_c_716_n 0.00585385f $X=1.87 $Y=2.465 $X2=0 $Y2=0
cc_264 N_B1_M1017_g N_VPWR_c_716_n 0.00486043f $X=2.3 $Y=2.465 $X2=0 $Y2=0
cc_265 N_B1_M1004_g N_VPWR_c_703_n 0.0108791f $X=1.87 $Y=2.465 $X2=0 $Y2=0
cc_266 N_B1_M1017_g N_VPWR_c_703_n 0.00458264f $X=2.3 $Y=2.465 $X2=0 $Y2=0
cc_267 N_B1_M1005_g N_A_32_65#_c_902_n 0.010819f $X=1.87 $Y=0.745 $X2=0 $Y2=0
cc_268 N_B1_M1015_g N_A_32_65#_c_902_n 0.0104125f $X=2.3 $Y=0.745 $X2=0 $Y2=0
cc_269 N_B1_c_287_n N_A_32_65#_c_902_n 0.0447809f $X=2.08 $Y=1.51 $X2=0 $Y2=0
cc_270 N_B1_c_288_n N_A_32_65#_c_902_n 0.00246333f $X=2.3 $Y=1.51 $X2=0 $Y2=0
cc_271 N_B1_M1005_g N_A_289_65#_c_948_n 0.00242267f $X=1.87 $Y=0.745 $X2=0 $Y2=0
cc_272 N_B1_M1005_g N_A_289_65#_c_953_n 0.0130206f $X=1.87 $Y=0.745 $X2=0 $Y2=0
cc_273 N_B1_M1015_g N_A_289_65#_c_953_n 0.00955132f $X=2.3 $Y=0.745 $X2=0 $Y2=0
cc_274 N_B1_M1015_g N_A_389_65#_c_970_n 0.00803088f $X=2.3 $Y=0.745 $X2=0 $Y2=0
cc_275 N_B1_M1005_g N_A_389_65#_c_974_n 0.00464897f $X=1.87 $Y=0.745 $X2=0 $Y2=0
cc_276 N_B1_M1015_g N_A_389_65#_c_974_n 0.0045696f $X=2.3 $Y=0.745 $X2=0 $Y2=0
cc_277 N_B1_M1005_g N_VGND_c_1041_n 0.00356225f $X=1.87 $Y=0.745 $X2=0 $Y2=0
cc_278 N_B1_M1015_g N_VGND_c_1041_n 0.00302901f $X=2.3 $Y=0.745 $X2=0 $Y2=0
cc_279 N_B1_M1005_g N_VGND_c_1049_n 0.00511014f $X=1.87 $Y=0.745 $X2=0 $Y2=0
cc_280 N_B1_M1015_g N_VGND_c_1049_n 0.00434735f $X=2.3 $Y=0.745 $X2=0 $Y2=0
cc_281 N_A2_M1006_g N_A1_c_454_n 0.0406753f $X=3.63 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A2_c_337_n N_A1_c_454_n 0.00608853f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_283 N_A2_c_342_n N_A1_c_454_n 0.0010862f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_284 A2 N_A1_c_454_n 5.71612e-19 $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_285 N_A2_c_338_n N_A1_c_455_n 0.0148511f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_286 N_A2_c_342_n N_A1_c_455_n 0.00612865f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A2_c_349_n N_A1_c_465_n 0.0328346f $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_288 N_A2_c_340_n N_A1_c_456_n 0.00699466f $X=4.995 $Y=1.65 $X2=0 $Y2=0
cc_289 N_A2_c_342_n N_A1_c_456_n 0.0087837f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A2_c_343_n N_A1_c_456_n 0.00175617f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A2_c_344_n N_A1_c_456_n 6.61908e-19 $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_292 N_A2_M1023_g N_A1_c_457_n 0.0212656f $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_293 N_A2_c_342_n N_A1_c_457_n 0.00612865f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A2_c_337_n N_A1_c_458_n 0.0110263f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_295 N_A2_c_342_n N_A1_c_458_n 0.0083718f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_296 A2 N_A1_c_458_n 8.28471e-19 $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_297 N_A2_c_340_n N_A1_c_459_n 0.00977434f $X=4.995 $Y=1.65 $X2=0 $Y2=0
cc_298 N_A2_M1006_g A1 0.00106898f $X=3.63 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A2_c_337_n A1 0.00207961f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_300 N_A2_c_340_n A1 0.00560292f $X=4.995 $Y=1.65 $X2=0 $Y2=0
cc_301 N_A2_c_342_n A1 0.0626795f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A2_c_343_n A1 0.00777683f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A2_c_344_n A1 8.09667e-19 $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_304 N_A2_c_345_n A1 9.85511e-19 $X=3.61 $Y=1.26 $X2=0 $Y2=0
cc_305 A2 A1 0.0295599f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_306 N_A2_M1006_g N_A1_c_461_n 8.02896e-19 $X=3.63 $Y=2.465 $X2=0 $Y2=0
cc_307 N_A2_c_343_n N_A1_c_461_n 6.30906e-19 $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A2_c_344_n N_A1_c_461_n 0.004261f $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_309 N_A2_c_345_n N_A1_c_461_n 0.00371131f $X=3.61 $Y=1.26 $X2=0 $Y2=0
cc_310 N_A2_M1023_g N_A_32_367#_M1003_g 0.0191933f $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_311 N_A2_c_343_n N_A_32_367#_M1003_g 0.00104501f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A2_c_344_n N_A_32_367#_M1002_g 0.00256078f $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_313 N_A2_M1006_g N_A_32_367#_c_581_n 0.0130017f $X=3.63 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A2_c_337_n N_A_32_367#_c_581_n 0.00353192f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_315 N_A2_c_349_n N_A_32_367#_c_581_n 0.0126581f $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_316 N_A2_c_345_n N_A_32_367#_c_581_n 2.01179e-19 $X=3.61 $Y=1.26 $X2=0 $Y2=0
cc_317 A2 N_A_32_367#_c_581_n 0.0148267f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_318 N_A2_c_349_n N_A_32_367#_c_537_n 2.73158e-19 $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_319 N_A2_c_343_n N_A_32_367#_c_537_n 0.0146009f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A2_c_344_n N_A_32_367#_c_537_n 0.00567127f $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_321 N_A2_c_349_n N_A_32_367#_c_525_n 5.87351e-19 $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_322 N_A2_c_344_n N_A_32_367#_c_525_n 0.00299663f $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_323 N_A2_c_343_n N_A_32_367#_c_526_n 0.0146075f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A2_c_344_n N_A_32_367#_c_526_n 6.92287e-19 $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_325 N_A2_c_345_n N_A_32_367#_c_573_n 3.73717e-19 $X=3.61 $Y=1.26 $X2=0 $Y2=0
cc_326 A2 N_A_32_367#_c_573_n 0.0133014f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_327 N_A2_c_349_n N_A_32_367#_c_540_n 0.00714524f $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_328 N_A2_c_339_n N_A_32_367#_c_540_n 0.00914578f $X=5.165 $Y=1.65 $X2=0 $Y2=0
cc_329 N_A2_c_342_n N_A_32_367#_c_540_n 0.00738583f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A2_c_343_n N_A_32_367#_c_540_n 0.0117019f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A2_c_343_n N_A_32_367#_c_527_n 8.27028e-19 $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A2_c_344_n N_A_32_367#_c_527_n 0.0217042f $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_333 N_A2_M1006_g N_VPWR_c_707_n 0.00122096f $X=3.63 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_c_349_n N_VPWR_c_707_n 0.00122096f $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_335 N_A2_c_349_n N_VPWR_c_708_n 0.0038257f $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_336 N_A2_M1006_g N_VPWR_c_712_n 0.00585385f $X=3.63 $Y=2.465 $X2=0 $Y2=0
cc_337 N_A2_c_349_n N_VPWR_c_717_n 0.00585385f $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_338 N_A2_M1006_g N_VPWR_c_703_n 0.0120903f $X=3.63 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A2_c_349_n N_VPWR_c_703_n 0.0120903f $X=4.92 $Y=1.725 $X2=0 $Y2=0
cc_340 N_A2_c_343_n N_X_c_840_n 0.0059797f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A2_c_345_n N_A_32_65#_c_902_n 2.96418e-19 $X=3.61 $Y=1.26 $X2=0 $Y2=0
cc_342 N_A2_c_346_n N_A_32_65#_c_902_n 0.0138496f $X=3.572 $Y=1.245 $X2=0 $Y2=0
cc_343 A2 N_A_32_65#_c_902_n 7.89834e-19 $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_344 N_A2_c_346_n N_A_32_65#_c_904_n 7.79017e-19 $X=3.572 $Y=1.245 $X2=0 $Y2=0
cc_345 N_A2_c_343_n N_A_389_65#_M1008_s 7.6787e-19 $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A2_c_338_n N_A_389_65#_c_971_n 0.00283046f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_347 N_A2_c_338_n N_A_389_65#_c_972_n 0.0124146f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_348 N_A2_c_342_n N_A_389_65#_c_972_n 0.0210563f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A2_c_345_n N_A_389_65#_c_972_n 0.00216329f $X=3.61 $Y=1.26 $X2=0 $Y2=0
cc_350 N_A2_c_346_n N_A_389_65#_c_972_n 0.0212732f $X=3.572 $Y=1.245 $X2=0 $Y2=0
cc_351 N_A2_c_345_n N_A_389_65#_c_973_n 4.46857e-19 $X=3.61 $Y=1.26 $X2=0 $Y2=0
cc_352 N_A2_c_346_n N_A_389_65#_c_973_n 0.0139988f $X=3.572 $Y=1.245 $X2=0 $Y2=0
cc_353 N_A2_c_342_n N_A_389_65#_c_989_n 0.0402255f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A2_M1023_g N_A_389_65#_c_990_n 0.00206864f $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_355 N_A2_c_342_n N_A_389_65#_c_990_n 0.0130216f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_356 N_A2_c_343_n N_A_389_65#_c_990_n 0.00562795f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_357 N_A2_c_344_n N_A_389_65#_c_990_n 2.08152e-19 $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_358 N_A2_M1023_g N_A_389_65#_c_994_n 0.00516273f $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_359 N_A2_c_342_n N_A_389_65#_c_995_n 0.0159074f $X=5.165 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A2_c_346_n N_VGND_M1019_s 0.00104255f $X=3.572 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_361 N_A2_c_338_n N_VGND_c_1034_n 0.00336413f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_362 N_A2_c_338_n N_VGND_c_1035_n 0.00437852f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_363 N_A2_c_338_n N_VGND_c_1036_n 5.51842e-19 $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_364 N_A2_M1023_g N_VGND_c_1036_n 4.78045e-19 $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_365 N_A2_M1023_g N_VGND_c_1037_n 0.00155098f $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_366 N_A2_c_343_n N_VGND_c_1037_n 0.00245861f $X=5.33 $Y=1.16 $X2=0 $Y2=0
cc_367 N_A2_c_344_n N_VGND_c_1037_n 4.04022e-19 $X=5.33 $Y=1.49 $X2=0 $Y2=0
cc_368 N_A2_M1023_g N_VGND_c_1043_n 0.0054895f $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_369 N_A2_c_338_n N_VGND_c_1049_n 0.00717581f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_370 N_A2_M1023_g N_VGND_c_1049_n 0.00991006f $X=5.31 $Y=0.655 $X2=0 $Y2=0
cc_371 N_A1_c_462_n N_A_32_367#_c_581_n 0.0104574f $X=4.06 $Y=1.725 $X2=0 $Y2=0
cc_372 N_A1_c_453_n N_A_32_367#_c_581_n 6.4135e-19 $X=4.305 $Y=1.65 $X2=0 $Y2=0
cc_373 N_A1_c_465_n N_A_32_367#_c_581_n 0.0105073f $X=4.49 $Y=1.725 $X2=0 $Y2=0
cc_374 N_A1_c_456_n N_A_32_367#_c_581_n 0.00166222f $X=4.805 $Y=1.26 $X2=0 $Y2=0
cc_375 N_A1_c_459_n N_A_32_367#_c_581_n 3.2597e-19 $X=4.47 $Y=1.65 $X2=0 $Y2=0
cc_376 A1 N_A_32_367#_c_581_n 0.0556921f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_377 N_A1_c_465_n N_A_32_367#_c_540_n 9.15296e-19 $X=4.49 $Y=1.725 $X2=0 $Y2=0
cc_378 N_A1_c_462_n N_VPWR_c_707_n 0.0119844f $X=4.06 $Y=1.725 $X2=0 $Y2=0
cc_379 N_A1_c_465_n N_VPWR_c_707_n 0.0119844f $X=4.49 $Y=1.725 $X2=0 $Y2=0
cc_380 N_A1_c_462_n N_VPWR_c_712_n 0.00486043f $X=4.06 $Y=1.725 $X2=0 $Y2=0
cc_381 N_A1_c_465_n N_VPWR_c_717_n 0.00486043f $X=4.49 $Y=1.725 $X2=0 $Y2=0
cc_382 N_A1_c_462_n N_VPWR_c_703_n 0.0082726f $X=4.06 $Y=1.725 $X2=0 $Y2=0
cc_383 N_A1_c_465_n N_VPWR_c_703_n 0.0082726f $X=4.49 $Y=1.725 $X2=0 $Y2=0
cc_384 N_A1_c_462_n N_A_741_367#_c_824_n 0.0122738f $X=4.06 $Y=1.725 $X2=0 $Y2=0
cc_385 N_A1_c_465_n N_A_741_367#_c_824_n 0.0122738f $X=4.49 $Y=1.725 $X2=0 $Y2=0
cc_386 N_A1_c_455_n N_A_389_65#_c_989_n 0.00990046f $X=4.45 $Y=1.185 $X2=0 $Y2=0
cc_387 N_A1_c_457_n N_A_389_65#_c_989_n 0.00986332f $X=4.88 $Y=1.185 $X2=0 $Y2=0
cc_388 N_A1_c_458_n N_A_389_65#_c_989_n 5.34223e-19 $X=4.47 $Y=1.26 $X2=0 $Y2=0
cc_389 N_A1_c_455_n N_VGND_c_1035_n 0.00365202f $X=4.45 $Y=1.185 $X2=0 $Y2=0
cc_390 N_A1_c_455_n N_VGND_c_1036_n 0.00772116f $X=4.45 $Y=1.185 $X2=0 $Y2=0
cc_391 N_A1_c_457_n N_VGND_c_1036_n 0.00779875f $X=4.88 $Y=1.185 $X2=0 $Y2=0
cc_392 N_A1_c_457_n N_VGND_c_1043_n 0.00365202f $X=4.88 $Y=1.185 $X2=0 $Y2=0
cc_393 N_A1_c_455_n N_VGND_c_1049_n 0.00434777f $X=4.45 $Y=1.185 $X2=0 $Y2=0
cc_394 N_A1_c_457_n N_VGND_c_1049_n 0.00434777f $X=4.88 $Y=1.185 $X2=0 $Y2=0
cc_395 N_A_32_367#_c_539_n N_VPWR_M1013_d 0.00176461f $X=1.145 $Y=1.98 $X2=-0.19
+ $Y2=-0.245
cc_396 N_A_32_367#_c_562_n N_VPWR_M1016_d 0.00516803f $X=1.945 $Y=2.375 $X2=0
+ $Y2=0
cc_397 N_A_32_367#_c_567_n N_VPWR_M1017_d 0.00350652f $X=2.85 $Y=2.38 $X2=0
+ $Y2=0
cc_398 N_A_32_367#_c_581_n N_VPWR_M1001_s 0.00336238f $X=4.97 $Y=2.015 $X2=0
+ $Y2=0
cc_399 N_A_32_367#_c_537_n N_VPWR_M1002_d 0.00270397f $X=5.675 $Y=1.84 $X2=0
+ $Y2=0
cc_400 N_A_32_367#_c_534_n N_VPWR_c_704_n 0.0170096f $X=0.56 $Y=1.9 $X2=0 $Y2=0
cc_401 N_A_32_367#_c_562_n N_VPWR_c_705_n 0.0200142f $X=1.945 $Y=2.375 $X2=0
+ $Y2=0
cc_402 N_A_32_367#_c_567_n N_VPWR_c_706_n 0.0167604f $X=2.85 $Y=2.38 $X2=0 $Y2=0
cc_403 N_A_32_367#_M1002_g N_VPWR_c_708_n 0.0152918f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_404 N_A_32_367#_M1009_g N_VPWR_c_708_n 7.24342e-19 $X=6.325 $Y=2.465 $X2=0
+ $Y2=0
cc_405 N_A_32_367#_c_536_n N_VPWR_c_708_n 0.0678608f $X=5.135 $Y=2.455 $X2=0
+ $Y2=0
cc_406 N_A_32_367#_c_537_n N_VPWR_c_708_n 0.0217948f $X=5.675 $Y=1.84 $X2=0
+ $Y2=0
cc_407 N_A_32_367#_c_527_n N_VPWR_c_708_n 3.91644e-19 $X=7.185 $Y=1.49 $X2=0
+ $Y2=0
cc_408 N_A_32_367#_M1002_g N_VPWR_c_709_n 7.27171e-19 $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_409 N_A_32_367#_M1009_g N_VPWR_c_709_n 0.0142791f $X=6.325 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_A_32_367#_M1014_g N_VPWR_c_709_n 0.0142791f $X=6.755 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A_32_367#_M1025_g N_VPWR_c_709_n 7.27171e-19 $X=7.185 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A_32_367#_M1014_g N_VPWR_c_711_n 7.27171e-19 $X=6.755 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A_32_367#_M1025_g N_VPWR_c_711_n 0.0153838f $X=7.185 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_A_32_367#_c_573_n N_VPWR_c_712_n 0.0468122f $X=3.197 $Y=2.38 $X2=0
+ $Y2=0
cc_415 N_A_32_367#_c_533_n N_VPWR_c_714_n 0.0178111f $X=0.285 $Y=2.91 $X2=0
+ $Y2=0
cc_416 N_A_32_367#_c_629_p N_VPWR_c_715_n 0.0136943f $X=1.145 $Y=2.465 $X2=0
+ $Y2=0
cc_417 N_A_32_367#_c_630_p N_VPWR_c_716_n 0.0140491f $X=2.085 $Y=2.91 $X2=0
+ $Y2=0
cc_418 N_A_32_367#_c_536_n N_VPWR_c_717_n 0.0188755f $X=5.135 $Y=2.455 $X2=0
+ $Y2=0
cc_419 N_A_32_367#_M1002_g N_VPWR_c_718_n 0.00486043f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_A_32_367#_M1009_g N_VPWR_c_718_n 0.00486043f $X=6.325 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_A_32_367#_M1014_g N_VPWR_c_719_n 0.00486043f $X=6.755 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_32_367#_M1025_g N_VPWR_c_719_n 0.00486043f $X=7.185 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_32_367#_M1013_s N_VPWR_c_703_n 0.00371702f $X=0.16 $Y=1.835 $X2=0
+ $Y2=0
cc_424 N_A_32_367#_M1026_s N_VPWR_c_703_n 0.0041489f $X=1.005 $Y=1.835 $X2=0
+ $Y2=0
cc_425 N_A_32_367#_M1004_s N_VPWR_c_703_n 0.00253254f $X=1.945 $Y=1.835 $X2=0
+ $Y2=0
cc_426 N_A_32_367#_M1022_s N_VPWR_c_703_n 0.00676438f $X=2.805 $Y=1.835 $X2=0
+ $Y2=0
cc_427 N_A_32_367#_M1024_s N_VPWR_c_703_n 0.0026734f $X=4.995 $Y=1.835 $X2=0
+ $Y2=0
cc_428 N_A_32_367#_M1002_g N_VPWR_c_703_n 0.00824727f $X=5.895 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A_32_367#_M1009_g N_VPWR_c_703_n 0.00824727f $X=6.325 $Y=2.465 $X2=0
+ $Y2=0
cc_430 N_A_32_367#_M1014_g N_VPWR_c_703_n 0.00824727f $X=6.755 $Y=2.465 $X2=0
+ $Y2=0
cc_431 N_A_32_367#_M1025_g N_VPWR_c_703_n 0.00824727f $X=7.185 $Y=2.465 $X2=0
+ $Y2=0
cc_432 N_A_32_367#_c_533_n N_VPWR_c_703_n 0.0100304f $X=0.285 $Y=2.91 $X2=0
+ $Y2=0
cc_433 N_A_32_367#_c_629_p N_VPWR_c_703_n 0.00866444f $X=1.145 $Y=2.465 $X2=0
+ $Y2=0
cc_434 N_A_32_367#_c_630_p N_VPWR_c_703_n 0.0090585f $X=2.085 $Y=2.91 $X2=0
+ $Y2=0
cc_435 N_A_32_367#_c_567_n N_VPWR_c_703_n 0.0107284f $X=2.85 $Y=2.38 $X2=0 $Y2=0
cc_436 N_A_32_367#_c_536_n N_VPWR_c_703_n 0.0111968f $X=5.135 $Y=2.455 $X2=0
+ $Y2=0
cc_437 N_A_32_367#_c_573_n N_VPWR_c_703_n 0.02702f $X=3.197 $Y=2.38 $X2=0 $Y2=0
cc_438 N_A_32_367#_c_581_n N_A_741_367#_M1006_d 0.00447479f $X=4.97 $Y=2.015
+ $X2=-0.19 $Y2=-0.245
cc_439 N_A_32_367#_c_581_n N_A_741_367#_M1011_d 0.00346223f $X=4.97 $Y=2.015
+ $X2=0 $Y2=0
cc_440 N_A_32_367#_c_581_n N_A_741_367#_c_824_n 0.0309139f $X=4.97 $Y=2.015
+ $X2=0 $Y2=0
cc_441 N_A_32_367#_c_581_n N_A_741_367#_c_829_n 0.0129403f $X=4.97 $Y=2.015
+ $X2=0 $Y2=0
cc_442 N_A_32_367#_c_581_n N_A_741_367#_c_830_n 0.0129403f $X=4.97 $Y=2.015
+ $X2=0 $Y2=0
cc_443 N_A_32_367#_M1010_g N_X_c_839_n 0.0138529f $X=6.21 $Y=0.655 $X2=0 $Y2=0
cc_444 N_A_32_367#_M1012_g N_X_c_839_n 0.014115f $X=6.64 $Y=0.655 $X2=0 $Y2=0
cc_445 N_A_32_367#_c_658_p N_X_c_839_n 0.0469271f $X=6.89 $Y=1.49 $X2=0 $Y2=0
cc_446 N_A_32_367#_c_527_n N_X_c_839_n 0.00289453f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_447 N_A_32_367#_M1003_g N_X_c_840_n 0.00252993f $X=5.78 $Y=0.655 $X2=0 $Y2=0
cc_448 N_A_32_367#_c_658_p N_X_c_840_n 0.0182231f $X=6.89 $Y=1.49 $X2=0 $Y2=0
cc_449 N_A_32_367#_c_527_n N_X_c_840_n 0.00299787f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_450 N_A_32_367#_M1009_g N_X_c_845_n 0.0130035f $X=6.325 $Y=2.465 $X2=0 $Y2=0
cc_451 N_A_32_367#_M1014_g N_X_c_845_n 0.0131657f $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_452 N_A_32_367#_c_658_p N_X_c_845_n 0.0598561f $X=6.89 $Y=1.49 $X2=0 $Y2=0
cc_453 N_A_32_367#_c_527_n N_X_c_845_n 0.00286055f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_454 N_A_32_367#_M1002_g N_X_c_846_n 6.54275e-19 $X=5.895 $Y=2.465 $X2=0 $Y2=0
cc_455 N_A_32_367#_c_537_n N_X_c_846_n 0.0106583f $X=5.675 $Y=1.84 $X2=0 $Y2=0
cc_456 N_A_32_367#_c_658_p N_X_c_846_n 0.0153881f $X=6.89 $Y=1.49 $X2=0 $Y2=0
cc_457 N_A_32_367#_c_527_n N_X_c_846_n 0.00296179f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_458 N_A_32_367#_M1020_g N_X_c_841_n 0.0168482f $X=7.07 $Y=0.655 $X2=0 $Y2=0
cc_459 N_A_32_367#_c_658_p N_X_c_841_n 0.00727995f $X=6.89 $Y=1.49 $X2=0 $Y2=0
cc_460 N_A_32_367#_c_527_n N_X_c_841_n 0.00297778f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_461 N_A_32_367#_c_658_p N_X_c_842_n 0.015388f $X=6.89 $Y=1.49 $X2=0 $Y2=0
cc_462 N_A_32_367#_c_527_n N_X_c_842_n 0.00299787f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_463 N_A_32_367#_M1025_g N_X_c_847_n 0.0155645f $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_464 N_A_32_367#_c_527_n N_X_c_847_n 0.00286055f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_465 N_A_32_367#_M1014_g X 4.82162e-19 $X=6.755 $Y=2.465 $X2=0 $Y2=0
cc_466 N_A_32_367#_M1020_g X 0.0036412f $X=7.07 $Y=0.655 $X2=0 $Y2=0
cc_467 N_A_32_367#_M1025_g X 0.00395244f $X=7.185 $Y=2.465 $X2=0 $Y2=0
cc_468 N_A_32_367#_c_658_p X 0.0136544f $X=6.89 $Y=1.49 $X2=0 $Y2=0
cc_469 N_A_32_367#_c_527_n X 0.0179385f $X=7.185 $Y=1.49 $X2=0 $Y2=0
cc_470 N_A_32_367#_M1018_s N_A_32_65#_c_900_n 0.00176461f $X=0.585 $Y=0.325
+ $X2=0 $Y2=0
cc_471 N_A_32_367#_c_535_n N_A_32_65#_c_900_n 0.0159805f $X=0.725 $Y=0.68 $X2=0
+ $Y2=0
cc_472 N_A_32_367#_c_573_n N_A_32_65#_c_902_n 0.00649382f $X=3.197 $Y=2.38 $X2=0
+ $Y2=0
cc_473 N_A_32_367#_c_535_n N_A_32_65#_c_903_n 0.0105582f $X=0.725 $Y=0.68 $X2=0
+ $Y2=0
cc_474 N_A_32_367#_c_539_n N_A_32_65#_c_903_n 0.00607789f $X=1.145 $Y=1.98 $X2=0
+ $Y2=0
cc_475 N_A_32_367#_M1003_g N_VGND_c_1037_n 0.00165353f $X=5.78 $Y=0.655 $X2=0
+ $Y2=0
cc_476 N_A_32_367#_M1003_g N_VGND_c_1038_n 6.45202e-19 $X=5.78 $Y=0.655 $X2=0
+ $Y2=0
cc_477 N_A_32_367#_M1010_g N_VGND_c_1038_n 0.0113454f $X=6.21 $Y=0.655 $X2=0
+ $Y2=0
cc_478 N_A_32_367#_M1012_g N_VGND_c_1038_n 0.0112648f $X=6.64 $Y=0.655 $X2=0
+ $Y2=0
cc_479 N_A_32_367#_M1020_g N_VGND_c_1038_n 6.30983e-19 $X=7.07 $Y=0.655 $X2=0
+ $Y2=0
cc_480 N_A_32_367#_M1012_g N_VGND_c_1040_n 6.30983e-19 $X=6.64 $Y=0.655 $X2=0
+ $Y2=0
cc_481 N_A_32_367#_M1020_g N_VGND_c_1040_n 0.0126581f $X=7.07 $Y=0.655 $X2=0
+ $Y2=0
cc_482 N_A_32_367#_M1003_g N_VGND_c_1044_n 0.00585385f $X=5.78 $Y=0.655 $X2=0
+ $Y2=0
cc_483 N_A_32_367#_M1010_g N_VGND_c_1044_n 0.00486043f $X=6.21 $Y=0.655 $X2=0
+ $Y2=0
cc_484 N_A_32_367#_M1012_g N_VGND_c_1045_n 0.00486043f $X=6.64 $Y=0.655 $X2=0
+ $Y2=0
cc_485 N_A_32_367#_M1020_g N_VGND_c_1045_n 0.00486043f $X=7.07 $Y=0.655 $X2=0
+ $Y2=0
cc_486 N_A_32_367#_M1003_g N_VGND_c_1049_n 0.0106414f $X=5.78 $Y=0.655 $X2=0
+ $Y2=0
cc_487 N_A_32_367#_M1010_g N_VGND_c_1049_n 0.00824727f $X=6.21 $Y=0.655 $X2=0
+ $Y2=0
cc_488 N_A_32_367#_M1012_g N_VGND_c_1049_n 0.00824727f $X=6.64 $Y=0.655 $X2=0
+ $Y2=0
cc_489 N_A_32_367#_M1020_g N_VGND_c_1049_n 0.00824727f $X=7.07 $Y=0.655 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_703_n N_A_741_367#_M1006_d 0.0041489f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_491 N_VPWR_c_703_n N_A_741_367#_M1011_d 0.00397496f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_M1001_s N_A_741_367#_c_824_n 0.00346959f $X=4.135 $Y=1.835 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_707_n N_A_741_367#_c_824_n 0.0170777f $X=4.275 $Y=2.745 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_712_n N_A_741_367#_c_829_n 0.0136943f $X=4.11 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_703_n N_A_741_367#_c_829_n 0.00866972f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_717_n N_A_741_367#_c_830_n 0.0138717f $X=5.515 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_703_n N_A_741_367#_c_830_n 0.00886411f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_703_n N_X_M1002_s 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_499 N_VPWR_c_703_n N_X_M1014_s 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_500 N_VPWR_c_718_n N_X_c_879_n 0.0124525f $X=6.375 $Y=3.33 $X2=0 $Y2=0
cc_501 N_VPWR_c_703_n N_X_c_879_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_502 N_VPWR_M1009_d N_X_c_845_n 0.00176461f $X=6.4 $Y=1.835 $X2=0 $Y2=0
cc_503 N_VPWR_c_709_n N_X_c_845_n 0.0170777f $X=6.54 $Y=2.18 $X2=0 $Y2=0
cc_504 N_VPWR_c_719_n N_X_c_883_n 0.0124525f $X=7.235 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_c_703_n N_X_c_883_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_M1025_d N_X_c_847_n 0.00262981f $X=7.26 $Y=1.835 $X2=0 $Y2=0
cc_507 N_VPWR_c_711_n N_X_c_847_n 0.0220026f $X=7.4 $Y=2.18 $X2=0 $Y2=0
cc_508 N_X_c_839_n N_VGND_M1010_d 0.00176461f $X=6.76 $Y=1.15 $X2=0 $Y2=0
cc_509 N_X_c_841_n N_VGND_M1020_d 3.40166e-19 $X=7.235 $Y=1.15 $X2=0 $Y2=0
cc_510 N_X_c_843_n N_VGND_M1020_d 0.00220592f $X=7.415 $Y=1.235 $X2=0 $Y2=0
cc_511 N_X_c_839_n N_VGND_c_1038_n 0.0170777f $X=6.76 $Y=1.15 $X2=0 $Y2=0
cc_512 N_X_c_841_n N_VGND_c_1040_n 0.00443444f $X=7.235 $Y=1.15 $X2=0 $Y2=0
cc_513 N_X_c_843_n N_VGND_c_1040_n 0.0193827f $X=7.415 $Y=1.235 $X2=0 $Y2=0
cc_514 N_X_c_893_p N_VGND_c_1044_n 0.0136943f $X=5.995 $Y=0.42 $X2=0 $Y2=0
cc_515 N_X_c_894_p N_VGND_c_1045_n 0.0124525f $X=6.855 $Y=0.42 $X2=0 $Y2=0
cc_516 N_X_M1003_s N_VGND_c_1049_n 0.0041489f $X=5.855 $Y=0.235 $X2=0 $Y2=0
cc_517 N_X_M1012_s N_VGND_c_1049_n 0.00536646f $X=6.715 $Y=0.235 $X2=0 $Y2=0
cc_518 N_X_c_893_p N_VGND_c_1049_n 0.00866972f $X=5.995 $Y=0.42 $X2=0 $Y2=0
cc_519 N_X_c_894_p N_VGND_c_1049_n 0.00730901f $X=6.855 $Y=0.42 $X2=0 $Y2=0
cc_520 N_A_32_65#_c_902_n N_A_289_65#_M1007_d 0.00250873f $X=2.85 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_521 N_A_32_65#_c_902_n N_A_289_65#_M1015_s 0.00176891f $X=2.85 $Y=1.17 $X2=0
+ $Y2=0
cc_522 N_A_32_65#_c_900_n N_A_289_65#_c_948_n 0.00709624f $X=1.06 $Y=0.34 $X2=0
+ $Y2=0
cc_523 N_A_32_65#_c_902_n N_A_289_65#_c_950_n 0.0209324f $X=2.85 $Y=1.17 $X2=0
+ $Y2=0
cc_524 N_A_32_65#_c_902_n N_A_289_65#_c_953_n 0.0466926f $X=2.85 $Y=1.17 $X2=0
+ $Y2=0
cc_525 N_A_32_65#_c_902_n N_A_389_65#_M1005_d 0.00176891f $X=2.85 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_526 N_A_32_65#_M1027_s N_A_389_65#_c_970_n 0.00428784f $X=2.805 $Y=0.325
+ $X2=0 $Y2=0
cc_527 N_A_32_65#_c_902_n N_A_389_65#_c_970_n 0.0027311f $X=2.85 $Y=1.17 $X2=0
+ $Y2=0
cc_528 N_A_32_65#_c_904_n N_A_389_65#_c_970_n 0.0240983f $X=3.015 $Y=0.7 $X2=0
+ $Y2=0
cc_529 N_A_32_65#_c_904_n N_A_389_65#_c_971_n 0.0102694f $X=3.015 $Y=0.7 $X2=0
+ $Y2=0
cc_530 N_A_32_65#_c_904_n N_A_389_65#_c_973_n 0.015923f $X=3.015 $Y=0.7 $X2=0
+ $Y2=0
cc_531 N_A_32_65#_c_900_n N_A_389_65#_c_974_n 8.81611e-19 $X=1.06 $Y=0.34 $X2=0
+ $Y2=0
cc_532 N_A_32_65#_c_900_n N_VGND_c_1041_n 0.0558492f $X=1.06 $Y=0.34 $X2=0 $Y2=0
cc_533 N_A_32_65#_c_901_n N_VGND_c_1041_n 0.0186386f $X=0.39 $Y=0.34 $X2=0 $Y2=0
cc_534 N_A_32_65#_c_900_n N_VGND_c_1049_n 0.0312041f $X=1.06 $Y=0.34 $X2=0 $Y2=0
cc_535 N_A_32_65#_c_901_n N_VGND_c_1049_n 0.0101082f $X=0.39 $Y=0.34 $X2=0 $Y2=0
cc_536 N_A_289_65#_c_953_n N_A_389_65#_M1005_d 0.00336039f $X=2.375 $Y=0.797
+ $X2=-0.19 $Y2=-0.245
cc_537 N_A_289_65#_M1015_s N_A_389_65#_c_970_n 0.00212094f $X=2.375 $Y=0.325
+ $X2=0 $Y2=0
cc_538 N_A_289_65#_c_951_n N_A_389_65#_c_970_n 0.00934397f $X=2.515 $Y=0.81
+ $X2=0 $Y2=0
cc_539 N_A_289_65#_c_953_n N_A_389_65#_c_970_n 0.00477839f $X=2.375 $Y=0.797
+ $X2=0 $Y2=0
cc_540 N_A_289_65#_c_948_n N_A_389_65#_c_974_n 0.0117536f $X=1.585 $Y=0.45 $X2=0
+ $Y2=0
cc_541 N_A_289_65#_c_953_n N_A_389_65#_c_974_n 0.0155435f $X=2.375 $Y=0.797
+ $X2=0 $Y2=0
cc_542 N_A_289_65#_c_948_n N_VGND_c_1041_n 0.0195642f $X=1.585 $Y=0.45 $X2=0
+ $Y2=0
cc_543 N_A_289_65#_c_953_n N_VGND_c_1041_n 0.00205823f $X=2.375 $Y=0.797 $X2=0
+ $Y2=0
cc_544 N_A_289_65#_c_948_n N_VGND_c_1049_n 0.012425f $X=1.585 $Y=0.45 $X2=0
+ $Y2=0
cc_545 N_A_289_65#_c_953_n N_VGND_c_1049_n 0.00479948f $X=2.375 $Y=0.797 $X2=0
+ $Y2=0
cc_546 N_A_389_65#_c_972_n N_VGND_M1019_s 0.00493947f $X=4.105 $Y=0.815
+ $X2=-0.19 $Y2=-0.245
cc_547 N_A_389_65#_c_989_n N_VGND_M1000_d 0.0032987f $X=5 $Y=0.82 $X2=0 $Y2=0
cc_548 N_A_389_65#_c_970_n N_VGND_c_1034_n 0.0144806f $X=3.35 $Y=0.34 $X2=0
+ $Y2=0
cc_549 N_A_389_65#_c_971_n N_VGND_c_1034_n 0.00908345f $X=3.435 $Y=0.725 $X2=0
+ $Y2=0
cc_550 N_A_389_65#_c_972_n N_VGND_c_1034_n 0.0147204f $X=4.105 $Y=0.815 $X2=0
+ $Y2=0
cc_551 N_A_389_65#_c_972_n N_VGND_c_1035_n 0.0021534f $X=4.105 $Y=0.815 $X2=0
+ $Y2=0
cc_552 N_A_389_65#_c_1018_p N_VGND_c_1035_n 0.0136557f $X=4.235 $Y=0.42 $X2=0
+ $Y2=0
cc_553 N_A_389_65#_c_989_n N_VGND_c_1035_n 0.00196209f $X=5 $Y=0.82 $X2=0 $Y2=0
cc_554 N_A_389_65#_c_989_n N_VGND_c_1036_n 0.016459f $X=5 $Y=0.82 $X2=0 $Y2=0
cc_555 N_A_389_65#_c_970_n N_VGND_c_1041_n 0.0821756f $X=3.35 $Y=0.34 $X2=0
+ $Y2=0
cc_556 N_A_389_65#_c_972_n N_VGND_c_1041_n 0.002573f $X=4.105 $Y=0.815 $X2=0
+ $Y2=0
cc_557 N_A_389_65#_c_974_n N_VGND_c_1041_n 0.0219872f $X=2.085 $Y=0.34 $X2=0
+ $Y2=0
cc_558 N_A_389_65#_c_989_n N_VGND_c_1043_n 0.00196209f $X=5 $Y=0.82 $X2=0 $Y2=0
cc_559 N_A_389_65#_c_994_n N_VGND_c_1043_n 0.0156443f $X=5.095 $Y=0.42 $X2=0
+ $Y2=0
cc_560 N_A_389_65#_M1019_d N_VGND_c_1049_n 0.00248633f $X=4.095 $Y=0.235 $X2=0
+ $Y2=0
cc_561 N_A_389_65#_M1008_s N_VGND_c_1049_n 0.00245017f $X=4.955 $Y=0.235 $X2=0
+ $Y2=0
cc_562 N_A_389_65#_c_970_n N_VGND_c_1049_n 0.0467035f $X=3.35 $Y=0.34 $X2=0
+ $Y2=0
cc_563 N_A_389_65#_c_972_n N_VGND_c_1049_n 0.00922589f $X=4.105 $Y=0.815 $X2=0
+ $Y2=0
cc_564 N_A_389_65#_c_1018_p N_VGND_c_1049_n 0.00865943f $X=4.235 $Y=0.42 $X2=0
+ $Y2=0
cc_565 N_A_389_65#_c_989_n N_VGND_c_1049_n 0.00891615f $X=5 $Y=0.82 $X2=0 $Y2=0
cc_566 N_A_389_65#_c_994_n N_VGND_c_1049_n 0.00983564f $X=5.095 $Y=0.42 $X2=0
+ $Y2=0
cc_567 N_A_389_65#_c_974_n N_VGND_c_1049_n 0.0122779f $X=2.085 $Y=0.34 $X2=0
+ $Y2=0
