* File: sky130_fd_sc_lp__o22ai_m.pxi.spice
* Created: Wed Sep  2 10:21:05 2020
* 
x_PM_SKY130_FD_SC_LP__O22AI_M%B1 N_B1_c_62_n N_B1_c_63_n N_B1_c_64_n N_B1_c_70_n
+ N_B1_c_71_n N_B1_c_65_n N_B1_M1004_g N_B1_M1001_g N_B1_c_66_n B1 B1 B1 B1 B1
+ B1 N_B1_c_68_n PM_SKY130_FD_SC_LP__O22AI_M%B1
x_PM_SKY130_FD_SC_LP__O22AI_M%B2 N_B2_M1006_g N_B2_M1002_g N_B2_c_106_n
+ N_B2_c_111_n B2 B2 B2 N_B2_c_108_n PM_SKY130_FD_SC_LP__O22AI_M%B2
x_PM_SKY130_FD_SC_LP__O22AI_M%A2 N_A2_M1007_g N_A2_M1000_g N_A2_c_149_n
+ N_A2_c_154_n A2 A2 A2 N_A2_c_151_n PM_SKY130_FD_SC_LP__O22AI_M%A2
x_PM_SKY130_FD_SC_LP__O22AI_M%A1 N_A1_M1005_g N_A1_M1003_g N_A1_c_198_n A1 A1 A1
+ A1 N_A1_c_196_n PM_SKY130_FD_SC_LP__O22AI_M%A1
x_PM_SKY130_FD_SC_LP__O22AI_M%VPWR N_VPWR_M1001_s N_VPWR_M1005_d N_VPWR_c_226_n
+ N_VPWR_c_227_n VPWR N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n
+ N_VPWR_c_225_n N_VPWR_c_232_n N_VPWR_c_233_n PM_SKY130_FD_SC_LP__O22AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O22AI_M%Y N_Y_M1004_d N_Y_M1002_d N_Y_c_268_n N_Y_c_269_n
+ N_Y_c_281_n N_Y_c_296_n N_Y_c_271_n N_Y_c_272_n Y
+ PM_SKY130_FD_SC_LP__O22AI_M%Y
x_PM_SKY130_FD_SC_LP__O22AI_M%A_85_82# N_A_85_82#_M1004_s N_A_85_82#_M1006_d
+ N_A_85_82#_M1003_d N_A_85_82#_c_324_n N_A_85_82#_c_333_n N_A_85_82#_c_325_n
+ N_A_85_82#_c_326_n N_A_85_82#_c_327_n N_A_85_82#_c_328_n
+ PM_SKY130_FD_SC_LP__O22AI_M%A_85_82#
x_PM_SKY130_FD_SC_LP__O22AI_M%VGND N_VGND_M1000_d N_VGND_c_359_n N_VGND_c_360_n
+ N_VGND_c_361_n VGND N_VGND_c_362_n N_VGND_c_363_n
+ PM_SKY130_FD_SC_LP__O22AI_M%VGND
cc_1 VNB N_B1_c_62_n 0.0031934f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.24
cc_2 VNB N_B1_c_63_n 0.0380201f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.015
cc_3 VNB N_B1_c_64_n 0.025141f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.015
cc_4 VNB N_B1_c_65_n 0.0182338f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.94
cc_5 VNB N_B1_c_66_n 0.0254181f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_6 VNB B1 0.0100537f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_B1_c_68_n 0.0380317f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_8 VNB N_B2_M1006_g 0.0386762f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.015
cc_9 VNB N_B2_c_106_n 0.0128633f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.885
cc_10 VNB B2 0.00192404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_c_108_n 0.018505f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_12 VNB N_A2_M1000_g 0.030511f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.94
cc_13 VNB N_A2_c_149_n 0.0197249f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.885
cc_14 VNB A2 0.00113197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_151_n 0.0166647f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_16 VNB N_A1_M1003_g 0.0629963f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.94
cc_17 VNB A1 0.019361f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_18 VNB N_A1_c_196_n 0.0110262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_225_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_20 VNB N_Y_c_268_n 0.00703202f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.94
cc_21 VNB N_Y_c_269_n 0.0116751f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.62
cc_22 VNB N_A_85_82#_c_324_n 0.00905766f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.39
cc_23 VNB N_A_85_82#_c_325_n 0.0230445f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_24 VNB N_A_85_82#_c_326_n 0.00722637f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_25 VNB N_A_85_82#_c_327_n 4.08405e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_26 VNB N_A_85_82#_c_328_n 0.019099f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.69
cc_27 VNB N_VGND_c_359_n 0.00659391f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=2.315
cc_28 VNB N_VGND_c_360_n 0.0494065f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.62
cc_29 VNB N_VGND_c_361_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.39
cc_30 VNB N_VGND_c_362_n 0.0232084f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_31 VNB N_VGND_c_363_n 0.201765f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.69
cc_32 VPB N_B1_c_62_n 0.0393723f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.24
cc_33 VPB N_B1_c_70_n 0.0475238f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.315
cc_34 VPB N_B1_c_71_n 0.0131151f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.315
cc_35 VPB N_B1_M1001_g 0.0286264f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.885
cc_36 VPB B1 0.0520858f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_37 VPB N_B2_M1002_g 0.0451846f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.94
cc_38 VPB N_B2_c_106_n 0.0144813f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.885
cc_39 VPB N_B2_c_111_n 0.0186935f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.885
cc_40 VPB B2 0.00192429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A2_M1007_g 0.0499184f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.015
cc_42 VPB N_A2_c_149_n 0.00417122f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.885
cc_43 VPB N_A2_c_154_n 0.0191015f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.885
cc_44 VPB A2 0.00654874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A1_M1005_g 0.0401334f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.015
cc_46 VPB N_A1_c_198_n 0.0728035f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.885
cc_47 VPB A1 0.0147524f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.61
cc_48 VPB N_A1_c_196_n 0.0107424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_226_n 0.0124195f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.62
cc_50 VPB N_VPWR_c_227_n 0.0128358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_228_n 0.0179462f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_52 VPB N_VPWR_c_229_n 0.0338385f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.69
cc_53 VPB N_VPWR_c_230_n 0.0159859f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.105
cc_54 VPB N_VPWR_c_225_n 0.069551f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.105
cc_55 VPB N_VPWR_c_232_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_233_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_57 VPB N_Y_c_269_n 0.0120932f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.62
cc_58 VPB N_Y_c_271_n 0.00237097f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.61
cc_59 VPB N_Y_c_272_n 0.0017184f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_60 VPB Y 0.00472851f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_61 N_B1_c_65_n N_B2_M1006_g 0.0223776f $X=0.845 $Y=0.94 $X2=0 $Y2=0
cc_62 N_B1_c_70_n N_B2_M1002_g 0.061466f $X=0.84 $Y=2.315 $X2=0 $Y2=0
cc_63 N_B1_c_66_n N_B2_c_106_n 0.002907f $X=0.27 $Y=1.61 $X2=0 $Y2=0
cc_64 N_B1_c_62_n N_B2_c_111_n 0.002907f $X=0.36 $Y=2.24 $X2=0 $Y2=0
cc_65 N_B1_c_68_n N_B2_c_108_n 0.002907f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B1_c_70_n N_VPWR_c_226_n 0.00665143f $X=0.84 $Y=2.315 $X2=0 $Y2=0
cc_67 N_B1_M1001_g N_VPWR_c_226_n 0.0102571f $X=0.915 $Y=2.885 $X2=0 $Y2=0
cc_68 B1 N_VPWR_c_226_n 0.00115588f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_69 B1 N_VPWR_c_228_n 0.0059365f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_B1_M1001_g N_VPWR_c_229_n 0.00486043f $X=0.915 $Y=2.885 $X2=0 $Y2=0
cc_71 N_B1_M1001_g N_VPWR_c_225_n 0.00445045f $X=0.915 $Y=2.885 $X2=0 $Y2=0
cc_72 B1 N_VPWR_c_225_n 0.00676397f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_B1_c_63_n N_Y_c_268_n 0.00385101f $X=0.77 $Y=1.015 $X2=0 $Y2=0
cc_74 N_B1_c_65_n N_Y_c_268_n 0.0155643f $X=0.845 $Y=0.94 $X2=0 $Y2=0
cc_75 B1 N_Y_c_268_n 0.00726911f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_B1_c_63_n N_Y_c_269_n 0.00814595f $X=0.77 $Y=1.015 $X2=0 $Y2=0
cc_77 N_B1_c_70_n N_Y_c_269_n 0.00809935f $X=0.84 $Y=2.315 $X2=0 $Y2=0
cc_78 B1 N_Y_c_269_n 0.0498805f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_79 N_B1_c_68_n N_Y_c_269_n 0.011689f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_80 N_B1_M1001_g N_Y_c_281_n 0.00404225f $X=0.915 $Y=2.885 $X2=0 $Y2=0
cc_81 N_B1_c_70_n N_Y_c_271_n 0.00415943f $X=0.84 $Y=2.315 $X2=0 $Y2=0
cc_82 N_B1_M1001_g N_Y_c_271_n 0.0044277f $X=0.915 $Y=2.885 $X2=0 $Y2=0
cc_83 B1 N_Y_c_271_n 0.00734011f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_B1_M1001_g N_Y_c_272_n 0.00469349f $X=0.915 $Y=2.885 $X2=0 $Y2=0
cc_85 N_B1_c_70_n Y 0.003671f $X=0.84 $Y=2.315 $X2=0 $Y2=0
cc_86 N_B1_M1001_g Y 0.00317468f $X=0.915 $Y=2.885 $X2=0 $Y2=0
cc_87 N_B1_c_65_n N_A_85_82#_c_324_n 0.0116881f $X=0.845 $Y=0.94 $X2=0 $Y2=0
cc_88 N_B1_c_64_n N_A_85_82#_c_328_n 0.0113482f $X=0.435 $Y=1.015 $X2=0 $Y2=0
cc_89 N_B1_c_65_n N_A_85_82#_c_328_n 0.00142375f $X=0.845 $Y=0.94 $X2=0 $Y2=0
cc_90 N_B1_c_65_n N_VGND_c_360_n 9.21892e-19 $X=0.845 $Y=0.94 $X2=0 $Y2=0
cc_91 B1 N_VGND_c_363_n 0.00780715f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_92 N_B2_c_111_n N_A2_M1007_g 0.0468776f $X=1.185 $Y=2 $X2=0 $Y2=0
cc_93 B2 N_A2_M1007_g 2.68982e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B2_M1006_g N_A2_M1000_g 0.0230274f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_95 N_B2_c_108_n N_A2_c_149_n 0.0115762f $X=1.185 $Y=1.495 $X2=0 $Y2=0
cc_96 N_B2_c_106_n N_A2_c_154_n 0.0115762f $X=1.185 $Y=1.835 $X2=0 $Y2=0
cc_97 N_B2_M1006_g A2 0.00248339f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_98 N_B2_c_111_n A2 0.00161317f $X=1.185 $Y=2 $X2=0 $Y2=0
cc_99 B2 A2 0.0403334f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B2_M1006_g N_A2_c_151_n 0.0115762f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_101 B2 N_A2_c_151_n 0.0022391f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B2_M1002_g N_VPWR_c_226_n 0.00205733f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_103 N_B2_M1002_g N_VPWR_c_229_n 0.00387146f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_104 N_B2_M1002_g N_VPWR_c_225_n 0.00540804f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_105 N_B2_M1006_g N_Y_c_268_n 0.00746284f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_106 B2 N_Y_c_268_n 0.00971283f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B2_c_108_n N_Y_c_268_n 0.00363823f $X=1.185 $Y=1.495 $X2=0 $Y2=0
cc_108 N_B2_M1006_g N_Y_c_269_n 0.00481078f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_109 N_B2_M1002_g N_Y_c_269_n 0.00476058f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_110 B2 N_Y_c_269_n 0.0635897f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B2_c_108_n N_Y_c_269_n 0.00746763f $X=1.185 $Y=1.495 $X2=0 $Y2=0
cc_112 N_B2_M1002_g N_Y_c_281_n 0.00375623f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_113 N_B2_M1002_g N_Y_c_296_n 0.00503229f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_114 N_B2_M1002_g N_Y_c_272_n 0.00571495f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_115 N_B2_M1002_g Y 0.00688921f $X=1.275 $Y=2.885 $X2=0 $Y2=0
cc_116 N_B2_c_111_n Y 0.0033945f $X=1.185 $Y=2 $X2=0 $Y2=0
cc_117 B2 Y 0.0142332f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B2_M1006_g N_A_85_82#_c_324_n 0.0140671f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_119 N_B2_M1006_g N_A_85_82#_c_333_n 0.0060828f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_120 N_B2_M1006_g N_A_85_82#_c_326_n 0.00158033f $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_121 N_B2_M1006_g N_VGND_c_360_n 9.21892e-19 $X=1.275 $Y=0.62 $X2=0 $Y2=0
cc_122 N_A2_M1000_g N_A1_M1003_g 0.0253676f $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_123 A2 N_A1_M1003_g 6.59882e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_124 N_A2_c_151_n N_A1_M1003_g 0.0116742f $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_125 N_A2_M1007_g N_A1_c_198_n 0.0774768f $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_126 N_A2_c_154_n N_A1_c_198_n 0.0116742f $X=1.755 $Y=1.88 $X2=0 $Y2=0
cc_127 A2 N_A1_c_198_n 7.56589e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A2_M1007_g A1 0.00286209f $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_129 A2 A1 0.0563707f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_151_n A1 0.00477283f $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_131 N_A2_c_149_n N_A1_c_196_n 0.0116742f $X=1.755 $Y=1.715 $X2=0 $Y2=0
cc_132 N_A2_M1007_g N_VPWR_c_227_n 0.0022041f $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_133 N_A2_M1007_g N_VPWR_c_229_n 0.00552362f $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_134 N_A2_M1007_g N_VPWR_c_225_n 0.00993496f $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_135 N_A2_M1000_g N_Y_c_268_n 2.03027e-19 $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_136 N_A2_M1007_g N_Y_c_296_n 0.00463555f $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_137 A2 N_Y_c_296_n 0.00133374f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A2_M1007_g N_Y_c_272_n 0.0011409f $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_139 N_A2_M1007_g Y 9.26079e-19 $X=1.705 $Y=2.885 $X2=0 $Y2=0
cc_140 N_A2_M1000_g N_A_85_82#_c_324_n 0.00125755f $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_141 N_A2_M1000_g N_A_85_82#_c_333_n 6.59275e-19 $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_142 N_A2_M1000_g N_A_85_82#_c_325_n 0.0123484f $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_143 A2 N_A_85_82#_c_325_n 0.0110607f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A2_c_151_n N_A_85_82#_c_325_n 0.00262118f $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_145 A2 N_A_85_82#_c_326_n 0.00622737f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A2_c_151_n N_A_85_82#_c_326_n 8.84835e-19 $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_147 N_A2_M1000_g N_VGND_c_359_n 0.00504771f $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_148 N_A2_M1000_g N_VGND_c_360_n 0.00529112f $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_149 N_A2_M1000_g N_VGND_c_363_n 0.00518865f $X=1.785 $Y=0.62 $X2=0 $Y2=0
cc_150 N_A1_M1005_g N_VPWR_c_227_n 0.0105915f $X=2.065 $Y=2.885 $X2=0 $Y2=0
cc_151 N_A1_c_198_n N_VPWR_c_227_n 0.00218418f $X=2.325 $Y=2.12 $X2=0 $Y2=0
cc_152 A1 N_VPWR_c_227_n 0.012128f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A1_M1005_g N_VPWR_c_229_n 0.00486043f $X=2.065 $Y=2.885 $X2=0 $Y2=0
cc_154 N_A1_M1005_g N_VPWR_c_225_n 0.0070005f $X=2.065 $Y=2.885 $X2=0 $Y2=0
cc_155 A1 N_VPWR_c_225_n 0.00284872f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A1_M1005_g N_Y_c_296_n 8.57853e-19 $X=2.065 $Y=2.885 $X2=0 $Y2=0
cc_157 N_A1_M1003_g N_A_85_82#_c_325_n 0.0131345f $X=2.235 $Y=0.62 $X2=0 $Y2=0
cc_158 A1 N_A_85_82#_c_325_n 0.0240456f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A1_c_196_n N_A_85_82#_c_325_n 0.00272742f $X=2.325 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_M1003_g N_A_85_82#_c_327_n 3.52891e-19 $X=2.235 $Y=0.62 $X2=0 $Y2=0
cc_161 N_A1_M1003_g N_VGND_c_359_n 0.0143839f $X=2.235 $Y=0.62 $X2=0 $Y2=0
cc_162 N_A1_M1003_g N_VGND_c_362_n 0.00455951f $X=2.235 $Y=0.62 $X2=0 $Y2=0
cc_163 N_A1_M1003_g N_VGND_c_363_n 0.00447788f $X=2.235 $Y=0.62 $X2=0 $Y2=0
cc_164 N_VPWR_c_225_n A_198_535# 0.00258157f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_165 N_VPWR_c_225_n N_Y_M1002_d 0.00246398f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VPWR_c_226_n N_Y_c_281_n 0.00482087f $X=0.7 $Y=2.95 $X2=0 $Y2=0
cc_167 N_VPWR_c_229_n N_Y_c_281_n 0.00487883f $X=2.115 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_225_n N_Y_c_281_n 0.00560863f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_169 N_VPWR_c_227_n N_Y_c_296_n 0.00275243f $X=2.28 $Y=2.95 $X2=0 $Y2=0
cc_170 N_VPWR_c_229_n N_Y_c_296_n 0.0103399f $X=2.115 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_225_n N_Y_c_296_n 0.0122047f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_226_n N_Y_c_271_n 0.00370167f $X=0.7 $Y=2.95 $X2=0 $Y2=0
cc_173 N_VPWR_c_225_n N_Y_c_271_n 0.00237734f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_c_225_n Y 0.00620929f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_175 N_VPWR_c_225_n A_356_535# 0.00899413f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_176 A_198_535# N_Y_c_281_n 0.00281311f $X=0.99 $Y=2.675 $X2=0.7 $Y2=2.95
cc_177 A_198_535# N_Y_c_272_n 4.40361e-19 $X=0.99 $Y=2.675 $X2=0.535 $Y2=3.33
cc_178 N_Y_M1004_d N_A_85_82#_c_324_n 0.00180746f $X=0.92 $Y=0.41 $X2=0 $Y2=0
cc_179 N_Y_c_268_n N_A_85_82#_c_324_n 0.0192361f $X=0.835 $Y=1.01 $X2=0 $Y2=0
cc_180 N_Y_c_268_n N_A_85_82#_c_333_n 0.0126904f $X=0.835 $Y=1.01 $X2=0 $Y2=0
cc_181 N_Y_c_268_n N_A_85_82#_c_326_n 0.0113949f $X=0.835 $Y=1.01 $X2=0 $Y2=0
cc_182 N_A_85_82#_c_324_n N_VGND_c_359_n 0.0123841f $X=1.465 $Y=0.355 $X2=0
+ $Y2=0
cc_183 N_A_85_82#_c_325_n N_VGND_c_359_n 0.0201653f $X=2.365 $Y=0.925 $X2=0
+ $Y2=0
cc_184 N_A_85_82#_c_324_n N_VGND_c_360_n 0.0579002f $X=1.465 $Y=0.355 $X2=0
+ $Y2=0
cc_185 N_A_85_82#_c_328_n N_VGND_c_360_n 0.0206108f $X=0.55 $Y=0.355 $X2=0 $Y2=0
cc_186 N_A_85_82#_c_327_n N_VGND_c_362_n 0.00463199f $X=2.45 $Y=0.685 $X2=0
+ $Y2=0
cc_187 N_A_85_82#_c_324_n N_VGND_c_363_n 0.0360461f $X=1.465 $Y=0.355 $X2=0
+ $Y2=0
cc_188 N_A_85_82#_c_325_n N_VGND_c_363_n 0.0126278f $X=2.365 $Y=0.925 $X2=0
+ $Y2=0
cc_189 N_A_85_82#_c_327_n N_VGND_c_363_n 0.00610964f $X=2.45 $Y=0.685 $X2=0
+ $Y2=0
cc_190 N_A_85_82#_c_328_n N_VGND_c_363_n 0.0124745f $X=0.55 $Y=0.355 $X2=0 $Y2=0
