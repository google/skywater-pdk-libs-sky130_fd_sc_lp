* NGSPICE file created from sky130_fd_sc_lp__a32o_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_432_47# B2 VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=1.1088e+12p ps=7.68e+06u
M1001 VGND a_108_267# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1002 a_631_47# A1 a_108_267# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=4.074e+11p ps=2.65e+06u
M1003 a_345_367# B1 a_108_267# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3923e+12p pd=9.77e+06u as=3.528e+11p ps=3.08e+06u
M1004 a_345_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.1592e+12p ps=9.4e+06u
M1005 VPWR a_108_267# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=6.678e+11p ps=6.1e+06u
M1006 X a_108_267# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_345_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_108_267# B2 a_345_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_739_47# A2 a_631_47# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1010 a_108_267# B1 a_432_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_108_267# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A3 a_345_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A3 a_739_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

