* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4_lp A B C D VGND VNB VPB VPWR X
X0 a_114_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_47# D a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND C a_272_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_154_419# C a_252_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_252_419# B a_366_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_366_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_27_47# A a_646_167# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_465_185# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_646_167# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_272_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_804_167# a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND B a_465_185# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_27_47# a_804_167# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_27_47# D a_154_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
