* File: sky130_fd_sc_lp__a221o_2.pxi.spice
* Created: Wed Sep  2 09:21:16 2020
* 
x_PM_SKY130_FD_SC_LP__A221O_2%A_86_27# N_A_86_27#_M1003_d N_A_86_27#_M1013_d
+ N_A_86_27#_M1010_s N_A_86_27#_c_73_n N_A_86_27#_M1011_g N_A_86_27#_M1004_g
+ N_A_86_27#_c_75_n N_A_86_27#_M1012_g N_A_86_27#_M1009_g N_A_86_27#_c_77_n
+ N_A_86_27#_c_78_n N_A_86_27#_c_79_n N_A_86_27#_c_147_p N_A_86_27#_c_80_n
+ N_A_86_27#_c_81_n N_A_86_27#_c_82_n N_A_86_27#_c_83_n N_A_86_27#_c_125_p
+ N_A_86_27#_c_87_n PM_SKY130_FD_SC_LP__A221O_2%A_86_27#
x_PM_SKY130_FD_SC_LP__A221O_2%A2 N_A2_c_174_n N_A2_M1000_g N_A2_M1008_g A2
+ N_A2_c_176_n PM_SKY130_FD_SC_LP__A221O_2%A2
x_PM_SKY130_FD_SC_LP__A221O_2%A1 N_A1_M1007_g N_A1_M1003_g A1 A1 N_A1_c_214_n
+ N_A1_c_217_n PM_SKY130_FD_SC_LP__A221O_2%A1
x_PM_SKY130_FD_SC_LP__A221O_2%C1 N_C1_M1013_g N_C1_M1010_g C1 N_C1_c_253_n
+ N_C1_c_256_n PM_SKY130_FD_SC_LP__A221O_2%C1
x_PM_SKY130_FD_SC_LP__A221O_2%B1 N_B1_M1006_g N_B1_M1005_g B1 N_B1_c_285_n
+ N_B1_c_286_n PM_SKY130_FD_SC_LP__A221O_2%B1
x_PM_SKY130_FD_SC_LP__A221O_2%B2 N_B2_M1001_g N_B2_M1002_g B2 B2 N_B2_c_322_n
+ N_B2_c_323_n PM_SKY130_FD_SC_LP__A221O_2%B2
x_PM_SKY130_FD_SC_LP__A221O_2%VPWR N_VPWR_M1004_s N_VPWR_M1009_s N_VPWR_M1007_d
+ N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n
+ VPWR N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_348_n N_VPWR_c_357_n
+ N_VPWR_c_358_n PM_SKY130_FD_SC_LP__A221O_2%VPWR
x_PM_SKY130_FD_SC_LP__A221O_2%X N_X_M1011_s N_X_M1004_d X X X X X X X
+ N_X_c_405_n PM_SKY130_FD_SC_LP__A221O_2%X
x_PM_SKY130_FD_SC_LP__A221O_2%A_334_367# N_A_334_367#_M1000_d
+ N_A_334_367#_M1005_d N_A_334_367#_c_424_n N_A_334_367#_c_423_n
+ N_A_334_367#_c_437_n N_A_334_367#_c_430_n
+ PM_SKY130_FD_SC_LP__A221O_2%A_334_367#
x_PM_SKY130_FD_SC_LP__A221O_2%A_653_367# N_A_653_367#_M1010_d
+ N_A_653_367#_M1002_d N_A_653_367#_c_458_n N_A_653_367#_c_456_n
+ N_A_653_367#_c_457_n PM_SKY130_FD_SC_LP__A221O_2%A_653_367#
x_PM_SKY130_FD_SC_LP__A221O_2%VGND N_VGND_M1011_d N_VGND_M1012_d N_VGND_M1013_s
+ N_VGND_M1001_d N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n
+ N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n VGND N_VGND_c_479_n
+ N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n
+ PM_SKY130_FD_SC_LP__A221O_2%VGND
cc_1 VNB N_A_86_27#_c_73_n 0.0213512f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.215
cc_2 VNB N_A_86_27#_M1004_g 0.00873618f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_3 VNB N_A_86_27#_c_75_n 0.0177815f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.215
cc_4 VNB N_A_86_27#_M1009_g 0.00625656f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_5 VNB N_A_86_27#_c_77_n 0.00538267f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.38
cc_6 VNB N_A_86_27#_c_78_n 0.0713314f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.38
cc_7 VNB N_A_86_27#_c_79_n 0.00949909f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.16
cc_8 VNB N_A_86_27#_c_80_n 0.0128529f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=0.42
cc_9 VNB N_A_86_27#_c_81_n 0.00893851f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=1.93
cc_10 VNB N_A_86_27#_c_82_n 0.0145652f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.165
cc_11 VNB N_A_86_27#_c_83_n 0.0226374f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.165
cc_12 VNB N_A2_c_174_n 0.0308298f $X=-0.19 $Y=-0.245 $X2=2.14 $Y2=0.265
cc_13 VNB N_A2_M1008_g 0.0180091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_176_n 0.00209376f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.545
cc_15 VNB N_A1_M1003_g 0.0264886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_214_n 0.0337475f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.215
cc_17 VNB N_C1_M1013_g 0.0276513f $X=-0.19 $Y=-0.245 $X2=2.85 $Y2=1.835
cc_18 VNB N_C1_c_253_n 0.0285661f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.685
cc_19 VNB N_B1_M1006_g 0.0243761f $X=-0.19 $Y=-0.245 $X2=2.85 $Y2=1.835
cc_20 VNB N_B1_c_285_n 0.0269218f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.685
cc_21 VNB N_B1_c_286_n 0.0017614f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.545
cc_22 VNB N_B2_M1002_g 0.0070637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B2 0.0327967f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.215
cc_24 VNB N_B2_c_322_n 0.0349722f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.215
cc_25 VNB N_B2_c_323_n 0.0218061f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.685
cc_26 VNB N_VPWR_c_348_n 0.203486f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=0.42
cc_27 VNB N_X_c_405_n 0.00539742f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_28 VNB N_VGND_c_472_n 0.0119587f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.545
cc_29 VNB N_VGND_c_473_n 0.0515715f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_30 VNB N_VGND_c_474_n 0.00276782f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.685
cc_31 VNB N_VGND_c_475_n 0.011339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_476_n 0.0342778f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.38
cc_33 VNB N_VGND_c_477_n 0.0272418f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.16
cc_34 VNB N_VGND_c_478_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.075
cc_35 VNB N_VGND_c_479_n 0.0148053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_480_n 0.032628f $X=-0.19 $Y=-0.245 $X2=3.44 $Y2=1.075
cc_37 VNB N_VGND_c_481_n 0.0126445f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.38
cc_38 VNB N_VGND_c_482_n 0.28826f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.38
cc_39 VNB N_VGND_c_483_n 0.0109159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_484_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A_86_27#_M1004_g 0.0272176f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_42 VPB N_A_86_27#_M1009_g 0.022375f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_43 VPB N_A_86_27#_c_81_n 0.00673821f $X=-0.19 $Y=1.655 $X2=2.67 $Y2=1.93
cc_44 VPB N_A_86_27#_c_87_n 0.00996953f $X=-0.19 $Y=1.655 $X2=2.975 $Y2=2.095
cc_45 VPB N_A2_c_174_n 0.00651729f $X=-0.19 $Y=1.655 $X2=2.14 $Y2=0.265
cc_46 VPB N_A2_M1000_g 0.021047f $X=-0.19 $Y=1.655 $X2=2.85 $Y2=1.835
cc_47 VPB N_A2_c_176_n 0.00578133f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.545
cc_48 VPB N_A1_M1007_g 0.0229511f $X=-0.19 $Y=1.655 $X2=2.85 $Y2=1.835
cc_49 VPB N_A1_c_214_n 0.00945895f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=1.215
cc_50 VPB N_A1_c_217_n 0.00557738f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.685
cc_51 VPB N_C1_M1010_g 0.0232379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_C1_c_253_n 0.00668913f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.685
cc_53 VPB N_C1_c_256_n 0.00273835f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.545
cc_54 VPB N_B1_M1005_g 0.0189607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B1_c_285_n 0.00635311f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.685
cc_56 VPB N_B1_c_286_n 0.00611935f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.545
cc_57 VPB N_B2_M1002_g 0.0262543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB B2 0.0159315f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.215
cc_59 VPB N_VPWR_c_349_n 0.0119328f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.215
cc_60 VPB N_VPWR_c_350_n 0.0666542f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.685
cc_61 VPB N_VPWR_c_351_n 0.00511587f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.685
cc_62 VPB N_VPWR_c_352_n 0.0168514f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_63 VPB N_VPWR_c_353_n 0.00751567f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.38
cc_64 VPB N_VPWR_c_354_n 0.0194732f $X=-0.19 $Y=1.655 $X2=1.235 $Y2=1.16
cc_65 VPB N_VPWR_c_355_n 0.0623717f $X=-0.19 $Y=1.655 $X2=3.44 $Y2=0.42
cc_66 VPB N_VPWR_c_348_n 0.0605542f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=0.42
cc_67 VPB N_VPWR_c_357_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.975 $Y2=2.095
cc_68 VPB N_VPWR_c_358_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.38
cc_69 VPB N_X_c_405_n 0.00415667f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_70 VPB N_A_334_367#_c_423_n 0.017697f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.545
cc_71 VPB N_A_653_367#_c_456_n 0.0131643f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.685
cc_72 VPB N_A_653_367#_c_457_n 0.0328646f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.545
cc_73 N_A_86_27#_M1009_g N_A2_c_174_n 0.00326359f $X=0.935 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_74 N_A_86_27#_c_77_n N_A2_c_174_n 0.00157021f $X=1.07 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_75 N_A_86_27#_c_78_n N_A2_c_174_n 0.0172097f $X=1.07 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_86_27#_c_79_n N_A2_c_174_n 0.00503021f $X=2.115 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A_86_27#_M1009_g N_A2_M1000_g 0.0261041f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_86_27#_c_75_n N_A2_M1008_g 0.00708003f $X=0.935 $Y=1.215 $X2=0 $Y2=0
cc_79 N_A_86_27#_c_78_n N_A2_M1008_g 8.38313e-19 $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_80 N_A_86_27#_c_79_n N_A2_M1008_g 0.0150149f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_86_27#_c_80_n N_A2_M1008_g 0.00261871f $X=2.28 $Y=0.42 $X2=0 $Y2=0
cc_82 N_A_86_27#_M1009_g N_A2_c_176_n 0.00115004f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_86_27#_c_77_n N_A2_c_176_n 0.00754489f $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_84 N_A_86_27#_c_78_n N_A2_c_176_n 4.8418e-19 $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_85 N_A_86_27#_c_79_n N_A2_c_176_n 0.027707f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_86_27#_c_81_n N_A1_M1007_g 9.9579e-19 $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_87 N_A_86_27#_c_87_n N_A1_M1007_g 0.00140951f $X=2.975 $Y=2.095 $X2=0 $Y2=0
cc_88 N_A_86_27#_c_79_n N_A1_M1003_g 0.0132888f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_86_27#_c_80_n N_A1_M1003_g 0.016683f $X=2.28 $Y=0.42 $X2=0 $Y2=0
cc_90 N_A_86_27#_c_81_n N_A1_M1003_g 0.00228024f $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_91 N_A_86_27#_c_83_n N_A1_M1003_g 0.00442573f $X=2.755 $Y=1.165 $X2=0 $Y2=0
cc_92 N_A_86_27#_c_79_n N_A1_c_214_n 2.23934e-19 $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_86_27#_c_81_n N_A1_c_214_n 0.00429855f $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_94 N_A_86_27#_c_83_n N_A1_c_214_n 0.0067887f $X=2.755 $Y=1.165 $X2=0 $Y2=0
cc_95 N_A_86_27#_c_79_n N_A1_c_217_n 0.00280444f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_86_27#_c_81_n N_A1_c_217_n 0.0374163f $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_97 N_A_86_27#_c_83_n N_A1_c_217_n 0.0245534f $X=2.755 $Y=1.165 $X2=0 $Y2=0
cc_98 N_A_86_27#_c_87_n N_A1_c_217_n 0.0271772f $X=2.975 $Y=2.095 $X2=0 $Y2=0
cc_99 N_A_86_27#_c_80_n N_C1_M1013_g 0.00409763f $X=2.28 $Y=0.42 $X2=0 $Y2=0
cc_100 N_A_86_27#_c_81_n N_C1_M1013_g 0.00248999f $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_101 N_A_86_27#_c_82_n N_C1_M1013_g 0.0166818f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_102 N_A_86_27#_c_81_n N_C1_M1010_g 0.00473364f $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_103 N_A_86_27#_c_81_n N_C1_c_253_n 0.00417225f $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_104 N_A_86_27#_c_82_n N_C1_c_253_n 0.00444593f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_105 N_A_86_27#_c_87_n N_C1_c_253_n 8.08174e-19 $X=2.975 $Y=2.095 $X2=0 $Y2=0
cc_106 N_A_86_27#_c_81_n N_C1_c_256_n 0.02447f $X=2.67 $Y=1.93 $X2=0 $Y2=0
cc_107 N_A_86_27#_c_82_n N_C1_c_256_n 0.0243464f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_108 N_A_86_27#_c_87_n N_C1_c_256_n 0.0109539f $X=2.975 $Y=2.095 $X2=0 $Y2=0
cc_109 N_A_86_27#_c_82_n N_B1_M1006_g 0.00581856f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_110 N_A_86_27#_c_125_p N_B1_M1006_g 0.0163995f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_111 N_A_86_27#_c_82_n N_B1_c_285_n 0.00179595f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_112 N_A_86_27#_c_82_n N_B1_c_286_n 0.0113914f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_113 N_A_86_27#_c_82_n B2 0.00196253f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_114 N_A_86_27#_c_82_n N_B2_c_323_n 6.51072e-19 $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_115 N_A_86_27#_c_125_p N_B2_c_323_n 0.00254502f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_116 N_A_86_27#_M1004_g N_VPWR_c_350_n 0.00929098f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_86_27#_M1009_g N_VPWR_c_351_n 0.0164006f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_86_27#_c_77_n N_VPWR_c_351_n 0.00590667f $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_119 N_A_86_27#_c_78_n N_VPWR_c_351_n 9.12831e-19 $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_120 N_A_86_27#_c_79_n N_VPWR_c_351_n 0.00599668f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_86_27#_M1004_g N_VPWR_c_354_n 0.00585385f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_86_27#_M1009_g N_VPWR_c_354_n 0.00585385f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_86_27#_M1010_s N_VPWR_c_348_n 0.00348066f $X=2.85 $Y=1.835 $X2=0
+ $Y2=0
cc_124 N_A_86_27#_M1004_g N_VPWR_c_348_n 0.0114685f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_86_27#_M1009_g N_VPWR_c_348_n 0.011381f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_86_27#_c_73_n N_X_c_405_n 0.00337465f $X=0.505 $Y=1.215 $X2=0 $Y2=0
cc_127 N_A_86_27#_M1004_g N_X_c_405_n 0.00795653f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_86_27#_c_75_n N_X_c_405_n 0.00159547f $X=0.935 $Y=1.215 $X2=0 $Y2=0
cc_129 N_A_86_27#_M1009_g N_X_c_405_n 0.00552732f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_86_27#_c_77_n N_X_c_405_n 0.0213301f $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_131 N_A_86_27#_c_78_n N_X_c_405_n 0.0293039f $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_132 N_A_86_27#_c_147_p N_X_c_405_n 0.0124645f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_86_27#_c_79_n N_A_334_367#_c_424_n 0.00211444f $X=2.115 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_86_27#_M1010_s N_A_334_367#_c_423_n 0.00701432f $X=2.85 $Y=1.835
+ $X2=0 $Y2=0
cc_135 N_A_86_27#_c_87_n N_A_334_367#_c_423_n 0.0368648f $X=2.975 $Y=2.095 $X2=0
+ $Y2=0
cc_136 N_A_86_27#_c_79_n N_VGND_M1012_d 0.00363856f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_86_27#_c_147_p N_VGND_M1012_d 0.00182736f $X=1.235 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_86_27#_c_82_n N_VGND_M1013_s 0.00225733f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_139 N_A_86_27#_c_73_n N_VGND_c_473_n 0.00710604f $X=0.505 $Y=1.215 $X2=0
+ $Y2=0
cc_140 N_A_86_27#_c_73_n N_VGND_c_474_n 5.92482e-19 $X=0.505 $Y=1.215 $X2=0
+ $Y2=0
cc_141 N_A_86_27#_c_75_n N_VGND_c_474_n 0.0115522f $X=0.935 $Y=1.215 $X2=0 $Y2=0
cc_142 N_A_86_27#_c_78_n N_VGND_c_474_n 0.0011364f $X=1.07 $Y=1.38 $X2=0 $Y2=0
cc_143 N_A_86_27#_c_79_n N_VGND_c_474_n 0.0292488f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_86_27#_c_147_p N_VGND_c_474_n 0.0166796f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_86_27#_c_80_n N_VGND_c_474_n 0.0229903f $X=2.28 $Y=0.42 $X2=0 $Y2=0
cc_146 N_A_86_27#_c_80_n N_VGND_c_475_n 0.0319169f $X=2.28 $Y=0.42 $X2=0 $Y2=0
cc_147 N_A_86_27#_c_82_n N_VGND_c_475_n 0.0220881f $X=3.31 $Y=1.165 $X2=0 $Y2=0
cc_148 N_A_86_27#_c_125_p N_VGND_c_476_n 0.0213555f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_149 N_A_86_27#_c_125_p N_VGND_c_477_n 0.015688f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_150 N_A_86_27#_c_73_n N_VGND_c_479_n 0.00555245f $X=0.505 $Y=1.215 $X2=0
+ $Y2=0
cc_151 N_A_86_27#_c_75_n N_VGND_c_479_n 0.00461019f $X=0.935 $Y=1.215 $X2=0
+ $Y2=0
cc_152 N_A_86_27#_c_80_n N_VGND_c_480_n 0.0234289f $X=2.28 $Y=0.42 $X2=0 $Y2=0
cc_153 N_A_86_27#_M1013_d N_VGND_c_482_n 0.00380103f $X=3.265 $Y=0.245 $X2=0
+ $Y2=0
cc_154 N_A_86_27#_c_73_n N_VGND_c_482_n 0.0112053f $X=0.505 $Y=1.215 $X2=0 $Y2=0
cc_155 N_A_86_27#_c_75_n N_VGND_c_482_n 0.00820187f $X=0.935 $Y=1.215 $X2=0
+ $Y2=0
cc_156 N_A_86_27#_c_80_n N_VGND_c_482_n 0.0126421f $X=2.28 $Y=0.42 $X2=0 $Y2=0
cc_157 N_A_86_27#_c_125_p N_VGND_c_482_n 0.00984745f $X=3.405 $Y=0.42 $X2=0
+ $Y2=0
cc_158 N_A_86_27#_c_79_n A_356_53# 0.00366293f $X=2.115 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A2_M1000_g N_A1_M1007_g 0.0156151f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_c_174_n N_A1_M1003_g 0.00351823f $X=1.595 $Y=1.675 $X2=0 $Y2=0
cc_161 N_A2_M1008_g N_A1_M1003_g 0.0693315f $X=1.705 $Y=0.685 $X2=0 $Y2=0
cc_162 N_A2_c_174_n N_A1_c_214_n 0.0219157f $X=1.595 $Y=1.675 $X2=0 $Y2=0
cc_163 N_A2_c_176_n N_A1_c_214_n 0.00236154f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A2_c_174_n N_A1_c_217_n 2.47447e-19 $X=1.595 $Y=1.675 $X2=0 $Y2=0
cc_165 N_A2_M1000_g N_A1_c_217_n 8.64502e-19 $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A2_c_176_n N_A1_c_217_n 0.0201276f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A2_M1000_g N_VPWR_c_351_n 0.0138365f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_M1000_g N_VPWR_c_352_n 0.0054895f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A2_M1000_g N_VPWR_c_353_n 4.84913e-19 $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_M1000_g N_VPWR_c_348_n 0.010609f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A2_c_176_n N_X_c_405_n 0.00612808f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A2_c_174_n N_A_334_367#_c_424_n 5.27063e-19 $X=1.595 $Y=1.675 $X2=0
+ $Y2=0
cc_173 N_A2_M1000_g N_A_334_367#_c_424_n 0.00663715f $X=1.595 $Y=2.465 $X2=0
+ $Y2=0
cc_174 N_A2_c_176_n N_A_334_367#_c_424_n 0.0135809f $X=1.61 $Y=1.51 $X2=0 $Y2=0
cc_175 N_A2_M1000_g N_A_334_367#_c_430_n 0.00754007f $X=1.595 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A2_M1008_g N_VGND_c_474_n 0.0162211f $X=1.705 $Y=0.685 $X2=0 $Y2=0
cc_177 N_A2_M1008_g N_VGND_c_480_n 0.00461019f $X=1.705 $Y=0.685 $X2=0 $Y2=0
cc_178 N_A2_M1008_g N_VGND_c_482_n 0.00806991f $X=1.705 $Y=0.685 $X2=0 $Y2=0
cc_179 N_A1_c_214_n N_C1_c_253_n 0.00520071f $X=2.24 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A1_c_217_n N_VPWR_M1007_d 0.00421288f $X=2.24 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A1_M1007_g N_VPWR_c_352_n 0.00364644f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A1_M1007_g N_VPWR_c_353_n 0.00810297f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A1_M1007_g N_VPWR_c_348_n 0.00441974f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A1_M1007_g N_A_334_367#_c_424_n 0.00477437f $X=2.06 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A1_c_217_n N_A_334_367#_c_424_n 0.0259155f $X=2.24 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A1_M1007_g N_A_334_367#_c_423_n 0.0147407f $X=2.06 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A1_c_217_n N_A_334_367#_c_423_n 0.0217548f $X=2.24 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A1_M1003_g N_VGND_c_474_n 0.0027902f $X=2.065 $Y=0.685 $X2=0 $Y2=0
cc_189 N_A1_M1003_g N_VGND_c_475_n 0.00317451f $X=2.065 $Y=0.685 $X2=0 $Y2=0
cc_190 N_A1_M1003_g N_VGND_c_480_n 0.00520505f $X=2.065 $Y=0.685 $X2=0 $Y2=0
cc_191 N_A1_M1003_g N_VGND_c_482_n 0.0107285f $X=2.065 $Y=0.685 $X2=0 $Y2=0
cc_192 N_C1_M1013_g N_B1_M1006_g 0.0239138f $X=3.19 $Y=0.665 $X2=0 $Y2=0
cc_193 N_C1_M1010_g N_B1_M1005_g 0.0528578f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_194 N_C1_c_253_n N_B1_c_285_n 0.0215729f $X=3.1 $Y=1.51 $X2=0 $Y2=0
cc_195 N_C1_c_256_n N_B1_c_285_n 2.88395e-19 $X=3.1 $Y=1.51 $X2=0 $Y2=0
cc_196 N_C1_c_253_n N_B1_c_286_n 0.00186964f $X=3.1 $Y=1.51 $X2=0 $Y2=0
cc_197 N_C1_c_256_n N_B1_c_286_n 0.0259188f $X=3.1 $Y=1.51 $X2=0 $Y2=0
cc_198 N_C1_M1010_g N_VPWR_c_353_n 0.0069181f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_199 N_C1_M1010_g N_VPWR_c_355_n 0.00425088f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_200 N_C1_M1010_g N_VPWR_c_348_n 0.00750519f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_201 N_C1_M1010_g N_A_334_367#_c_423_n 0.0161877f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_202 N_C1_c_256_n N_A_334_367#_c_423_n 0.00395317f $X=3.1 $Y=1.51 $X2=0 $Y2=0
cc_203 N_C1_M1010_g N_A_334_367#_c_437_n 0.00187381f $X=3.19 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_C1_M1010_g N_A_653_367#_c_458_n 0.0148075f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_205 N_C1_M1013_g N_VGND_c_475_n 0.0137419f $X=3.19 $Y=0.665 $X2=0 $Y2=0
cc_206 N_C1_M1013_g N_VGND_c_477_n 0.00477554f $X=3.19 $Y=0.665 $X2=0 $Y2=0
cc_207 N_C1_M1013_g N_VGND_c_482_n 0.00828349f $X=3.19 $Y=0.665 $X2=0 $Y2=0
cc_208 N_B1_M1005_g N_B2_M1002_g 0.0311564f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B1_c_286_n N_B2_M1002_g 2.67445e-19 $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_210 N_B1_M1006_g B2 0.00247583f $X=3.62 $Y=0.665 $X2=0 $Y2=0
cc_211 N_B1_M1005_g B2 2.40806e-19 $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_212 N_B1_c_285_n B2 0.00362218f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_213 N_B1_c_286_n B2 0.0255488f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_214 N_B1_c_285_n N_B2_c_322_n 0.0206187f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_215 N_B1_c_286_n N_B2_c_322_n 3.0266e-19 $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_216 N_B1_M1006_g N_B2_c_323_n 0.0446446f $X=3.62 $Y=0.665 $X2=0 $Y2=0
cc_217 N_B1_M1005_g N_VPWR_c_355_n 0.00357877f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B1_M1005_g N_VPWR_c_348_n 0.00553653f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B1_M1005_g N_A_334_367#_c_423_n 0.0118084f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B1_M1005_g N_A_334_367#_c_437_n 0.00978334f $X=3.62 $Y=2.465 $X2=0
+ $Y2=0
cc_221 N_B1_c_285_n N_A_334_367#_c_437_n 5.59281e-19 $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_222 N_B1_c_286_n N_A_334_367#_c_437_n 0.00879552f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_223 N_B1_M1005_g N_A_653_367#_c_458_n 0.0115665f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B1_M1006_g N_VGND_c_475_n 0.00127263f $X=3.62 $Y=0.665 $X2=0 $Y2=0
cc_225 N_B1_M1006_g N_VGND_c_476_n 0.00337427f $X=3.62 $Y=0.665 $X2=0 $Y2=0
cc_226 N_B1_M1006_g N_VGND_c_477_n 0.00539298f $X=3.62 $Y=0.665 $X2=0 $Y2=0
cc_227 N_B1_M1006_g N_VGND_c_482_n 0.0101168f $X=3.62 $Y=0.665 $X2=0 $Y2=0
cc_228 N_B2_M1002_g N_VPWR_c_355_n 0.00357877f $X=4.09 $Y=2.465 $X2=0 $Y2=0
cc_229 N_B2_M1002_g N_VPWR_c_348_n 0.00657127f $X=4.09 $Y=2.465 $X2=0 $Y2=0
cc_230 N_B2_M1002_g N_A_653_367#_c_458_n 0.0165264f $X=4.09 $Y=2.465 $X2=0 $Y2=0
cc_231 B2 N_A_653_367#_c_457_n 0.0245763f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_232 N_B2_c_322_n N_A_653_367#_c_457_n 7.27731e-19 $X=4.18 $Y=1.36 $X2=0 $Y2=0
cc_233 B2 N_VGND_c_476_n 0.0260007f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_234 N_B2_c_322_n N_VGND_c_476_n 0.0040906f $X=4.18 $Y=1.36 $X2=0 $Y2=0
cc_235 N_B2_c_323_n N_VGND_c_476_n 0.0239813f $X=4.18 $Y=1.195 $X2=0 $Y2=0
cc_236 N_B2_c_323_n N_VGND_c_477_n 0.00477554f $X=4.18 $Y=1.195 $X2=0 $Y2=0
cc_237 N_B2_c_323_n N_VGND_c_482_n 0.00842334f $X=4.18 $Y=1.195 $X2=0 $Y2=0
cc_238 N_VPWR_c_348_n N_X_M1004_d 0.00432284f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_350_n N_X_c_405_n 0.00152254f $X=0.29 $Y=1.98 $X2=0 $Y2=0
cc_240 N_VPWR_c_354_n N_X_c_405_n 0.0135169f $X=1.105 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_c_348_n N_X_c_405_n 0.00847534f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_348_n N_A_334_367#_M1000_d 0.00272835f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_243 N_VPWR_c_348_n N_A_334_367#_M1005_d 0.00257355f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_351_n N_A_334_367#_c_424_n 0.0330402f $X=1.27 $Y=2.005 $X2=0
+ $Y2=0
cc_245 N_VPWR_M1007_d N_A_334_367#_c_423_n 0.00552554f $X=2.135 $Y=1.835 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_352_n N_A_334_367#_c_423_n 0.00198381f $X=2.11 $Y=3.33 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_353_n N_A_334_367#_c_423_n 0.01532f $X=2.275 $Y=2.95 $X2=0 $Y2=0
cc_248 N_VPWR_c_355_n N_A_334_367#_c_423_n 0.0112309f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_348_n N_A_334_367#_c_423_n 0.0266394f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_351_n N_A_334_367#_c_430_n 0.0429461f $X=1.27 $Y=2.005 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_352_n N_A_334_367#_c_430_n 0.0181427f $X=2.11 $Y=3.33 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_348_n N_A_334_367#_c_430_n 0.0112063f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_348_n N_A_653_367#_M1010_d 0.00223577f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_254 N_VPWR_c_348_n N_A_653_367#_M1002_d 0.00211942f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_355_n N_A_653_367#_c_458_n 0.0534582f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_348_n N_A_653_367#_c_458_n 0.033719f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_355_n N_A_653_367#_c_456_n 0.0193375f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_348_n N_A_653_367#_c_456_n 0.0116633f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_X_c_405_n N_VGND_c_473_n 0.00224375f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_260 N_X_c_405_n N_VGND_c_474_n 0.0275297f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_261 N_X_c_405_n N_VGND_c_479_n 0.0156277f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_262 N_X_c_405_n N_VGND_c_482_n 0.00847534f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_263 N_A_334_367#_c_423_n N_A_653_367#_M1010_d 0.00805965f $X=3.67 $Y=2.515
+ $X2=-0.19 $Y2=1.655
cc_264 N_A_334_367#_M1005_d N_A_653_367#_c_458_n 0.00419917f $X=3.695 $Y=1.835
+ $X2=0 $Y2=0
cc_265 N_A_334_367#_c_423_n N_A_653_367#_c_458_n 0.040917f $X=3.67 $Y=2.515
+ $X2=0 $Y2=0
cc_266 N_VGND_c_482_n A_739_49# 0.0137053f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
