* File: sky130_fd_sc_lp__a2bb2o_1.pex.spice
* Created: Fri Aug 28 09:55:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%A_91_269# 1 2 9 13 16 17 18 19 21 23 26 29
+ 31 36
r96 36 38 11.1619 $w=2.83e-07 $l=2.3e-07 $layer=LI1_cond $X=2.592 $Y=0.445
+ $X2=2.592 $Y2=0.675
r97 33 34 14.1373 $w=2.33e-07 $l=2.7e-07 $layer=LI1_cond $X=2.217 $Y=2.14
+ $X2=2.217 $Y2=2.41
r98 29 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.62 $Y=1.51
+ $X2=0.62 $Y2=1.675
r99 29 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.62 $Y=1.51
+ $X2=0.62 $Y2=1.345
r100 28 31 8.45125 $w=2.98e-07 $l=2.2e-07 $layer=LI1_cond $X=0.62 $Y=1.495
+ $X2=0.84 $Y2=1.495
r101 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.51 $X2=0.62 $Y2=1.51
r102 26 38 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.65 $Y=2.055
+ $X2=2.65 $Y2=0.675
r103 24 33 2.58477 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.365 $Y=2.14
+ $X2=2.217 $Y2=2.14
r104 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.565 $Y=2.14
+ $X2=2.65 $Y2=2.055
r105 23 24 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.565 $Y=2.14
+ $X2=2.365 $Y2=2.14
r106 19 34 4.08828 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.217 $Y=2.495
+ $X2=2.217 $Y2=2.41
r107 19 21 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=2.217 $Y=2.495
+ $X2=2.217 $Y2=2.855
r108 17 34 2.58477 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.07 $Y=2.41
+ $X2=2.217 $Y2=2.41
r109 17 18 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=2.07 $Y=2.41
+ $X2=0.925 $Y2=2.41
r110 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.84 $Y=2.325
+ $X2=0.925 $Y2=2.41
r111 15 31 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.84 $Y=1.645 $X2=0.84
+ $Y2=1.495
r112 15 16 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.84 $Y=1.645
+ $X2=0.84 $Y2=2.325
r113 13 41 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.685 $Y=2.465
+ $X2=0.685 $Y2=1.675
r114 9 40 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.59 $Y=0.655
+ $X2=0.59 $Y2=1.345
r115 2 21 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=2.645 $X2=2.235 $Y2=2.855
r116 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.565 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%A1_N 2 5 9 11 12 13 14 15 16 23
r48 23 25 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.197 $Y=1.17
+ $X2=1.197 $Y2=1.005
r49 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.205
+ $Y=1.17 $X2=1.205 $Y2=1.17
r50 15 16 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.2
+ $Y2=2.035
r51 14 15 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r52 14 24 7.29665 $w=1.88e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=1.295
+ $X2=1.2 $Y2=1.17
r53 13 24 14.3014 $w=1.88e-07 $l=2.45e-07 $layer=LI1_cond $X=1.2 $Y=0.925
+ $X2=1.2 $Y2=1.17
r54 12 13 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.555 $X2=1.2
+ $Y2=0.925
r55 9 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.28 $Y=2.045
+ $X2=1.28 $Y2=1.675
r56 5 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.28 $Y=0.445
+ $X2=1.28 $Y2=1.005
r57 2 11 45.1798 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=1.197 $Y=1.503
+ $X2=1.197 $Y2=1.675
r58 1 23 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=1.197 $Y=1.177
+ $X2=1.197 $Y2=1.17
r59 1 2 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=1.197 $Y=1.177
+ $X2=1.197 $Y2=1.503
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%A2_N 3 7 11 12 13 16 17
r49 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.76 $Y=1.1
+ $X2=1.76 $Y2=1.1
r50 13 17 1.8762 $w=5.08e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.27 $X2=1.76
+ $Y2=1.27
r51 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.76 $Y=1.44
+ $X2=1.76 $Y2=1.1
r52 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.44
+ $X2=1.76 $Y2=1.605
r53 10 16 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=0.935
+ $X2=1.76 $Y2=1.1
r54 7 10 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.765 $Y=0.445
+ $X2=1.765 $Y2=0.935
r55 3 12 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.67 $Y=2.045
+ $X2=1.67 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%A_271_47# 1 2 9 15 19 20 21 22 25 27 28 31
+ 34 35 37 39
c90 39 0 1.47006e-19 $X=2.247 $Y=1.005
c91 37 0 1.46768e-19 $X=1.885 $Y=1.98
c92 27 0 1.45411e-19 $X=2.11 $Y=0.75
c93 25 0 6.51563e-20 $X=1.55 $Y=0.445
c94 22 0 6.54297e-20 $X=2.42 $Y=2.29
r95 37 38 16.7924 $w=2.63e-07 $l=3.62e-07 $layer=LI1_cond $X=1.885 $Y=1.875
+ $X2=2.247 $Y2=1.875
r96 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.3 $Y=1.17
+ $X2=2.3 $Y2=1.17
r97 32 38 0.46577 $w=2.75e-07 $l=1.7e-07 $layer=LI1_cond $X=2.247 $Y=1.705
+ $X2=2.247 $Y2=1.875
r98 32 34 22.4203 $w=2.73e-07 $l=5.35e-07 $layer=LI1_cond $X=2.247 $Y=1.705
+ $X2=2.247 $Y2=1.17
r99 31 39 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.247 $Y=1.142
+ $X2=2.247 $Y2=1.005
r100 31 34 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=2.247 $Y=1.142
+ $X2=2.247 $Y2=1.17
r101 29 39 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.195 $Y=0.835
+ $X2=2.195 $Y2=1.005
r102 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=0.75
+ $X2=2.195 $Y2=0.835
r103 27 28 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.11 $Y=0.75
+ $X2=1.715 $Y2=0.75
r104 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.59 $Y=0.665
+ $X2=1.715 $Y2=0.75
r105 23 25 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=1.59 $Y=0.665
+ $X2=1.59 $Y2=0.445
r106 21 22 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=2.42 $Y=2.14
+ $X2=2.42 $Y2=2.29
r107 20 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.39 $Y=1.675
+ $X2=2.39 $Y2=2.14
r108 19 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.3 $Y=1.51 $X2=2.3
+ $Y2=1.17
r109 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.51
+ $X2=2.3 $Y2=1.675
r110 18 35 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.005
+ $X2=2.3 $Y2=1.17
r111 15 22 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.45 $Y=2.855
+ $X2=2.45 $Y2=2.29
r112 9 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.35 $Y=0.445
+ $X2=2.35 $Y2=1.005
r113 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=1.835 $X2=1.885 $Y2=1.98
r114 1 25 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=1.355
+ $Y=0.235 $X2=1.55 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%B2 3 7 9 10 11 12 13 20
c49 20 0 1.46768e-19 $X=3 $Y=1.395
c50 9 0 6.54297e-20 $X=3.12 $Y=0.555
c51 3 0 2.92417e-19 $X=2.78 $Y=0.445
r52 20 23 88.3231 $w=4.6e-07 $l=5.05e-07 $layer=POLY_cond $X=2.935 $Y=1.395
+ $X2=2.935 $Y2=1.9
r53 20 22 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.935 $Y=1.395
+ $X2=2.935 $Y2=1.23
r54 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3 $Y=1.395
+ $X2=3 $Y2=1.395
r55 12 13 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.065 $Y=1.665
+ $X2=3.065 $Y2=2.035
r56 12 21 10.372 $w=2.98e-07 $l=2.7e-07 $layer=LI1_cond $X=3.065 $Y=1.665
+ $X2=3.065 $Y2=1.395
r57 11 21 3.84148 $w=2.98e-07 $l=1e-07 $layer=LI1_cond $X=3.065 $Y=1.295
+ $X2=3.065 $Y2=1.395
r58 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.065 $Y=0.925
+ $X2=3.065 $Y2=1.295
r59 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.065 $Y=0.555
+ $X2=3.065 $Y2=0.925
r60 7 23 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=2.88 $Y=2.855
+ $X2=2.88 $Y2=1.9
r61 3 22 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.78 $Y=0.445
+ $X2=2.78 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%B1 3 7 9 10 12 15 19 20 21 22 23 29
r40 22 23 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=2.035
r41 21 22 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.665
r42 20 21 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=0.925
+ $X2=3.57 $Y2=1.295
r43 20 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.005 $X2=3.57 $Y2=1.005
r44 18 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.005
r45 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.345
+ $X2=3.57 $Y2=1.51
r46 17 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.57 $Y=0.99
+ $X2=3.57 $Y2=1.005
r47 13 15 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.31 $Y=2.185
+ $X2=3.48 $Y2=2.185
r48 12 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.48 $Y=2.11
+ $X2=3.48 $Y2=2.185
r49 12 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.48 $Y=2.11 $X2=3.48
+ $Y2=1.51
r50 9 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.405 $Y=0.915
+ $X2=3.57 $Y2=0.99
r51 9 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=3.405 $Y=0.915
+ $X2=3.245 $Y2=0.915
r52 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.31 $Y=2.26 $X2=3.31
+ $Y2=2.185
r53 5 7 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=3.31 $Y=2.26 $X2=3.31
+ $Y2=2.855
r54 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.17 $Y=0.84
+ $X2=3.245 $Y2=0.915
r55 1 3 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.17 $Y=0.84 $X2=3.17
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%X 1 2 11 14 15 16 17 23 29
r25 21 29 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=0.305 $Y=0.895
+ $X2=0.305 $Y2=0.925
r26 17 31 7.65015 $w=3.98e-07 $l=1.43e-07 $layer=LI1_cond $X=0.305 $Y=0.952
+ $X2=0.305 $Y2=1.095
r27 17 29 0.777899 $w=3.98e-07 $l=2.7e-08 $layer=LI1_cond $X=0.305 $Y=0.952
+ $X2=0.305 $Y2=0.925
r28 17 21 0.80671 $w=3.98e-07 $l=2.8e-08 $layer=LI1_cond $X=0.305 $Y=0.867
+ $X2=0.305 $Y2=0.895
r29 16 17 8.98906 $w=3.98e-07 $l=3.12e-07 $layer=LI1_cond $X=0.305 $Y=0.555
+ $X2=0.305 $Y2=0.867
r30 16 23 3.8895 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=0.305 $Y=0.555
+ $X2=0.305 $Y2=0.42
r31 15 31 44.3636 $w=1.78e-07 $l=7.2e-07 $layer=LI1_cond $X=0.195 $Y=1.815
+ $X2=0.195 $Y2=1.095
r32 14 15 8.88815 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.335 $Y=1.98
+ $X2=0.335 $Y2=1.815
r33 9 14 1.69011 $w=4.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.335 $Y=2.045
+ $X2=0.335 $Y2=1.98
r34 9 11 22.4915 $w=4.58e-07 $l=8.65e-07 $layer=LI1_cond $X=0.335 $Y=2.045
+ $X2=0.335 $Y2=2.91
r35 2 14 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.835 $X2=0.47 $Y2=1.98
r36 2 11 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.835 $X2=0.47 $Y2=2.91
r37 1 23 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.25
+ $Y=0.235 $X2=0.375 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%VPWR 1 2 9 13 16 17 18 24 33 34 37
r40 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 34 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 31 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.095 $Y2=3.33
r44 31 33 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.26 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=3.095 $Y2=3.33
r50 24 29 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 18 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 16 21 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.9 $Y2=3.33
r57 15 26 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.9 $Y2=3.33
r59 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.095 $Y2=3.33
r60 11 13 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.095 $Y2=2.855
r61 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=3.245 $X2=0.9
+ $Y2=3.33
r62 7 9 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.9 $Y=3.245 $X2=0.9
+ $Y2=2.79
r63 2 13 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=2.645 $X2=3.095 $Y2=2.855
r64 1 9 600 $w=1.7e-07 $l=1.02261e-06 $layer=licon1_PDIFF $count=1 $X=0.76
+ $Y=1.835 $X2=0.9 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%A_505_529# 1 2 9 11 12 15
r25 13 15 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.56 $Y=2.565
+ $X2=3.56 $Y2=2.855
r26 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.43 $Y=2.48
+ $X2=3.56 $Y2=2.565
r27 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.43 $Y=2.48
+ $X2=2.76 $Y2=2.48
r28 7 12 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=2.647 $Y=2.565
+ $X2=2.76 $Y2=2.48
r29 7 9 14.8537 $w=2.23e-07 $l=2.9e-07 $layer=LI1_cond $X=2.647 $Y=2.565
+ $X2=2.647 $Y2=2.855
r30 2 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=2.645 $X2=3.525 $Y2=2.855
r31 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=2.645 $X2=2.665 $Y2=2.855
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_1%VGND 1 2 3 14 20 22 24 26 28 33 39 42 46
r57 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r59 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r60 37 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r61 37 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r62 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 34 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.055
+ $Y2=0
r64 34 36 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=3.12
+ $Y2=0
r65 33 45 4.09313 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.612
+ $Y2=0
r66 33 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.12
+ $Y2=0
r67 32 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r68 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 29 39 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.805
+ $Y2=0
r70 29 31 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.68
+ $Y2=0
r71 28 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.055
+ $Y2=0
r72 28 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r73 26 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r74 26 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r75 22 45 3.19156 $w=2.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.612 $Y2=0
r76 22 24 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.52 $Y2=0.445
r77 18 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r78 18 20 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.395
r79 14 16 24.3786 $w=2.58e-07 $l=5.5e-07 $layer=LI1_cond $X=0.805 $Y=0.38
+ $X2=0.805 $Y2=0.93
r80 12 39 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0
r81 12 14 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0.38
r82 3 24 182 $w=1.7e-07 $l=3.33879e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.49 $Y2=0.445
r83 2 20 182 $w=1.7e-07 $l=2.83945e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=2.055 $Y2=0.395
r84 1 16 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=0.665
+ $Y=0.235 $X2=0.805 $Y2=0.93
r85 1 14 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.665
+ $Y=0.235 $X2=0.805 $Y2=0.38
.ends

