* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4b_4 A_N B C D VGND VNB VPB VPWR X
X0 VPWR B a_242_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND a_242_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_825_49# a_49_133# a_242_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_242_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_242_23# a_49_133# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 X a_242_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND a_242_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 X a_242_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND D a_645_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_49_133# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR D a_242_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_645_49# C a_717_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_717_49# B a_825_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_49_133# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 X a_242_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR a_242_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VPWR a_242_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_242_23# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
