* File: sky130_fd_sc_lp__dlrtp_lp.spice
* Created: Fri Aug 28 10:27:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dlrtp_lp  VNB VPB GATE D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1010 A_114_57# N_GATE_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_186_57#_M1001_d N_GATE_M1001_g A_114_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_408_73# N_A_186_57#_M1006_g N_A_294_547#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.2086 PD=0.63 PS=1.92 NRD=14.28 NRS=34.284 M=1 R=2.8
+ SA=75000.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_186_57#_M1002_g A_408_73# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1019 A_566_73# N_D_M1019_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1020 N_A_638_73#_M1020_d N_D_M1020_g A_566_73# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_A_887_343#_M1028_d N_A_186_57#_M1028_g N_A_862_101#_M1028_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.168 PD=0.7 PS=1.64 NRD=0 NRS=32.856 M=1 R=2.8
+ SA=75000.3 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1026 A_1058_101# N_A_294_547#_M1026_g N_A_887_343#_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_638_73#_M1014_g A_1058_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1029 N_A_862_101#_M1029_d N_A_1208_75#_M1029_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_1510_47# N_A_887_343#_M1015_g N_A_1208_75#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1008 AS=0.2394 PD=1.08 PS=2.25 NRD=9.276 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1021 N_VGND_M1021_d N_RESET_B_M1021_g A_1510_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.5019 AS=0.1008 PD=2.035 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1016 A_1857_47# N_A_1208_75#_M1016_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.5019 PD=1.05 PS=2.035 NRD=7.14 NRS=130.704 M=1 R=5.6 SA=75001.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1007 N_Q_M1007_d N_A_1208_75#_M1007_g A_1857_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.0882 PD=2.3 PS=1.05 NRD=3.564 NRS=7.14 M=1 R=5.6 SA=75002.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 A_114_470# N_GATE_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1018 N_A_186_57#_M1018_d N_GATE_M1018_g A_114_470# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 A_384_345# N_A_186_57#_M1004_g N_A_294_547#_M1004_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=38.4741 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_186_57#_M1005_g A_384_345# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1616 AS=0.1152 PD=1.145 PS=1 NRD=0 NRS=38.4741 M=1 R=4.26667 SA=75000.7
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1008 A_617_345# N_D_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1616 PD=0.85 PS=1.145 NRD=15.3857 NRS=69.2455 M=1 R=4.26667 SA=75001.4
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_638_73#_M1011_d N_D_M1011_g A_617_345# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.7
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_887_343#_M1017_d N_A_186_57#_M1017_g N_A_800_343#_M1017_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.138023 AS=0.1824 PD=1.24981 PS=1.85 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1027 N_A_996_343#_M1027_d N_A_294_547#_M1027_g N_A_887_343#_M1017_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1197 AS=0.0905774 PD=1.41 PS=0.820189 NRD=0
+ NRS=53.9386 M=1 R=2.8 SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_638_73#_M1000_g N_A_800_343#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.138023 AS=0.1824 PD=1.24981 PS=1.85 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_996_343#_M1009_d N_A_1208_75#_M1009_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0905774 PD=1.41 PS=0.820189 NRD=0 NRS=56.2829 M=1
+ R=2.8 SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_887_343#_M1025_g N_A_1420_367#_M1025_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.4 A=0.189 P=2.82 MULT=1
MM1012 A_1593_367# N_RESET_B_M1012_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001 A=0.189 P=2.82 MULT=1
MM1013 N_A_1208_75#_M1013_d N_RESET_B_M1013_g A_1593_367# VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_A_1420_367#_M1003_d N_A_887_343#_M1003_g N_A_1208_75#_M1013_d VPB
+ PHIGHVT L=0.15 W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1
+ R=8.4 SA=75001.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1023 A_1949_367# N_A_1208_75#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3591 PD=1.5 PS=3.09 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1024 N_Q_M1024_d N_A_1208_75#_M1024_g A_1949_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1512 PD=3.09 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX30_noxref VNB VPB NWDIODE A=20.8747 P=25.85
c_165 VPB 0 1.43074e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlrtp_lp.pxi.spice"
*
.ends
*
*
