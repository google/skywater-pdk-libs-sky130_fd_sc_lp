* File: sky130_fd_sc_lp__a2111oi_2.spice
* Created: Wed Sep  2 09:16:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111oi_2.pex.spice"
.subckt sky130_fd_sc_lp__a2111oi_2  VNB VPB C1 D1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* D1	D1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1012 N_Y_M1012_d N_C1_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.7 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1012_s N_D1_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.2 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_D1_M1015_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1176 PD=1.23 PS=1.12 NRD=7.848 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003.8 A=0.126 P=1.98 MULT=1
MM1017 N_Y_M1017_d N_C1_M1017_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1365 AS=0.1638 PD=1.165 PS=1.23 NRD=4.284 NRS=7.848 M=1 R=5.6 SA=75001.6
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1017_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1365 PD=1.23 PS=1.165 NRD=5.712 NRS=2.136 M=1 R=5.6 SA=75002.1
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1003_d N_B1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1176 PD=1.23 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_684_47#_M1000_d N_A1_M1000_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.231 AS=0.1176 PD=1.39 PS=1.12 NRD=19.284 NRS=0 M=1 R=5.6 SA=75003
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1004 N_A_684_47#_M1000_d N_A2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.231 AS=0.1449 PD=1.39 PS=1.185 NRD=19.284 NRS=4.284 M=1 R=5.6 SA=75003.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1019 N_A_684_47#_M1019_d N_A2_M1019_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1449 PD=1.12 PS=1.185 NRD=0 NRS=4.992 M=1 R=5.6 SA=75004.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1013 N_A_684_47#_M1019_d N_A1_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75004.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_32_367#_M1005_d N_C1_M1005_g N_A_115_367#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1009 N_A_115_367#_M1005_s N_D1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1016 N_A_115_367#_M1016_d N_D1_M1016_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_A_32_367#_M1008_d N_C1_M1008_g N_A_115_367#_M1016_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1001 N_A_467_367#_M1001_d N_B1_M1001_g N_A_32_367#_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=6.2449 M=1 R=8.4 SA=75002
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_467_367#_M1001_d N_B1_M1010_g N_A_32_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_467_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_A_467_367#_M1006_d N_A2_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1018 N_A_467_367#_M1006_d N_A2_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1018_s N_A1_M1014_g N_A_467_367#_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.3339 PD=1.58 PS=3.05 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__a2111oi_2.pxi.spice"
*
.ends
*
*
