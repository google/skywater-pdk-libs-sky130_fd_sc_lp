* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2oi_lp A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR B2 a_27_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_494_47# A2_N a_296_146# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_296_146# A1_N a_652_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_652_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_409# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VGND A2_N a_494_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_409# a_296_146# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_456_339# A2_N a_296_146# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_456_339# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_170_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 Y a_296_146# a_334_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND B1 a_170_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_334_47# a_296_146# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
