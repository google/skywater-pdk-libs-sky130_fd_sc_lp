* File: sky130_fd_sc_lp__mux2_1.pxi.spice
* Created: Fri Aug 28 10:43:41 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_1%A_105_22# N_A_105_22#_M1001_d N_A_105_22#_M1005_d
+ N_A_105_22#_M1002_g N_A_105_22#_M1006_g N_A_105_22#_c_71_n N_A_105_22#_c_72_n
+ N_A_105_22#_c_73_n N_A_105_22#_c_117_p N_A_105_22#_c_74_n N_A_105_22#_c_75_n
+ N_A_105_22#_c_76_n PM_SKY130_FD_SC_LP__MUX2_1%A_105_22#
x_PM_SKY130_FD_SC_LP__MUX2_1%S N_S_M1007_g N_S_M1004_g N_S_M1003_g N_S_M1011_g
+ N_S_c_137_n N_S_c_144_n N_S_c_138_n N_S_c_139_n N_S_c_146_n N_S_c_147_n
+ N_S_c_148_n N_S_c_149_n S N_S_c_150_n N_S_c_151_n S
+ PM_SKY130_FD_SC_LP__MUX2_1%S
x_PM_SKY130_FD_SC_LP__MUX2_1%A1 N_A1_M1001_g N_A1_M1009_g N_A1_c_230_n
+ N_A1_c_231_n A1 A1 A1 A1 A1 A1 N_A1_c_232_n N_A1_c_236_n N_A1_c_233_n A1
+ PM_SKY130_FD_SC_LP__MUX2_1%A1
x_PM_SKY130_FD_SC_LP__MUX2_1%A0 N_A0_M1005_g N_A0_M1010_g A0 A0 A0 N_A0_c_294_n
+ PM_SKY130_FD_SC_LP__MUX2_1%A0
x_PM_SKY130_FD_SC_LP__MUX2_1%A_488_106# N_A_488_106#_M1003_d
+ N_A_488_106#_M1011_d N_A_488_106#_M1008_g N_A_488_106#_c_332_n
+ N_A_488_106#_c_333_n N_A_488_106#_M1000_g N_A_488_106#_c_335_n
+ N_A_488_106#_c_341_n N_A_488_106#_c_336_n N_A_488_106#_c_337_n
+ N_A_488_106#_c_338_n N_A_488_106#_c_339_n
+ PM_SKY130_FD_SC_LP__MUX2_1%A_488_106#
x_PM_SKY130_FD_SC_LP__MUX2_1%X N_X_M1002_s N_X_M1006_s X X X X X X X N_X_c_389_n
+ PM_SKY130_FD_SC_LP__MUX2_1%X
x_PM_SKY130_FD_SC_LP__MUX2_1%VPWR N_VPWR_M1006_d N_VPWR_M1000_d N_VPWR_c_402_n
+ N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n VPWR N_VPWR_c_406_n
+ N_VPWR_c_401_n N_VPWR_c_408_n PM_SKY130_FD_SC_LP__MUX2_1%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_1%VGND N_VGND_M1002_d N_VGND_M1008_d N_VGND_c_443_n
+ N_VGND_c_444_n VGND N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n
+ N_VGND_c_448_n N_VGND_c_449_n PM_SKY130_FD_SC_LP__MUX2_1%VGND
cc_1 VNB N_A_105_22#_M1006_g 0.0082546f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_2 VNB N_A_105_22#_c_71_n 0.00391395f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.355
cc_3 VNB N_A_105_22#_c_72_n 0.0396097f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.355
cc_4 VNB N_A_105_22#_c_73_n 0.0112622f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.075
cc_5 VNB N_A_105_22#_c_74_n 0.0115167f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=2.375
cc_6 VNB N_A_105_22#_c_75_n 0.00365759f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.87
cc_7 VNB N_A_105_22#_c_76_n 0.0213175f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.19
cc_8 VNB N_S_M1007_g 0.0303975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_S_M1003_g 0.0533138f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_10 VNB N_S_c_137_n 0.0122286f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.075
cc_11 VNB N_S_c_138_n 2.77691e-19 $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=2.375
cc_12 VNB N_S_c_139_n 0.0183479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_230_n 0.0183055f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.66
cc_14 VNB N_A1_c_231_n 0.0464562f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_15 VNB N_A1_c_232_n 0.0158224f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.355
cc_16 VNB N_A1_c_233_n 0.00559752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A1 0.0104378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A0_M1010_g 0.0385126f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.19
cc_19 VNB A0 0.00541516f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.66
cc_20 VNB N_A0_c_294_n 0.0180303f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.075
cc_21 VNB N_A_488_106#_M1008_g 0.0204389f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.66
cc_22 VNB N_A_488_106#_c_332_n 0.0310483f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_23 VNB N_A_488_106#_c_333_n 0.00724238f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_24 VNB N_A_488_106#_M1000_g 0.0064898f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.355
cc_25 VNB N_A_488_106#_c_335_n 0.00660126f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=1.355
cc_26 VNB N_A_488_106#_c_336_n 0.023597f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.355
cc_27 VNB N_A_488_106#_c_337_n 0.005391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_488_106#_c_338_n 0.0309436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_488_106#_c_339_n 0.0327026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_389_n 0.0716434f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=2.375
cc_31 VNB N_VPWR_c_401_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_443_n 0.00839109f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_33 VNB N_VGND_c_444_n 0.0331199f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.355
cc_34 VNB N_VGND_c_445_n 0.0497643f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.075
cc_35 VNB N_VGND_c_446_n 0.0268389f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.19
cc_36 VNB N_VGND_c_447_n 0.277414f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.52
cc_37 VNB N_VGND_c_448_n 0.0233828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_449_n 0.0113485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_105_22#_M1006_g 0.0270313f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_40 VPB N_A_105_22#_c_74_n 0.00539937f $X=-0.19 $Y=1.655 $X2=2.185 $Y2=2.375
cc_41 VPB N_S_M1004_g 0.0198008f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.19
cc_42 VPB N_S_M1003_g 0.00154742f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_43 VPB N_S_M1011_g 0.0260756f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.355
cc_44 VPB N_S_c_137_n 0.0144596f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.075
cc_45 VPB N_S_c_144_n 0.0197921f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.075
cc_46 VPB N_S_c_138_n 0.00891108f $X=-0.19 $Y=1.655 $X2=2.185 $Y2=2.375
cc_47 VPB N_S_c_146_n 0.0543982f $X=-0.19 $Y=1.655 $X2=1.94 $Y2=0.87
cc_48 VPB N_S_c_147_n 0.00351031f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=1.16
cc_49 VPB N_S_c_148_n 0.00354185f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.355
cc_50 VPB N_S_c_149_n 0.00869064f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.19
cc_51 VPB N_S_c_150_n 0.0361756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_S_c_151_n 0.0174087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A1_M1009_g 0.0224903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A1_c_236_n 0.0348735f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.52
cc_55 VPB A1 0.00305405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A0_M1005_g 0.0246674f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB A0 0.00496969f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=0.66
cc_58 VPB N_A0_c_294_n 0.0374836f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.075
cc_59 VPB N_A_488_106#_M1000_g 0.0364191f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.355
cc_60 VPB N_A_488_106#_c_341_n 0.0206717f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=2.375
cc_61 VPB N_A_488_106#_c_337_n 0.0312945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_X_c_389_n 0.0674439f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=2.375
cc_63 VPB N_VPWR_c_402_n 0.0190904f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_64 VPB N_VPWR_c_403_n 0.0286075f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.075
cc_65 VPB N_VPWR_c_404_n 0.0537063f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=2.375
cc_66 VPB N_VPWR_c_405_n 0.0043981f $X=-0.19 $Y=1.655 $X2=2.185 $Y2=2.375
cc_67 VPB N_VPWR_c_406_n 0.0270918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_401_n 0.0863769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_408_n 0.0270707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 N_A_105_22#_c_71_n N_S_M1007_g 0.00156934f $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_71 N_A_105_22#_c_72_n N_S_M1007_g 0.0072089f $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_72 N_A_105_22#_c_73_n N_S_M1007_g 0.0161864f $X=1.775 $Y=1.075 $X2=0 $Y2=0
cc_73 N_A_105_22#_c_75_n N_S_M1007_g 0.00136799f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_74 N_A_105_22#_c_76_n N_S_M1007_g 0.00933093f $X=0.712 $Y=1.19 $X2=0 $Y2=0
cc_75 N_A_105_22#_M1006_g N_S_M1004_g 0.00731395f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A_105_22#_M1006_g N_S_c_137_n 0.0097715f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_105_22#_M1006_g N_S_c_138_n 0.00148977f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_105_22#_c_71_n N_S_c_138_n 0.00820685f $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_79 N_A_105_22#_c_72_n N_S_c_138_n 5.70577e-19 $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_80 N_A_105_22#_c_73_n N_S_c_138_n 0.0123302f $X=1.775 $Y=1.075 $X2=0 $Y2=0
cc_81 N_A_105_22#_c_71_n N_S_c_139_n 6.63628e-19 $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_82 N_A_105_22#_c_72_n N_S_c_139_n 0.0112105f $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_83 N_A_105_22#_c_73_n N_S_c_139_n 0.00637215f $X=1.775 $Y=1.075 $X2=0 $Y2=0
cc_84 N_A_105_22#_c_74_n N_S_c_139_n 0.00235944f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_85 N_A_105_22#_c_74_n N_S_c_146_n 0.00940796f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_86 N_A_105_22#_c_73_n N_A1_c_230_n 0.00669296f $X=1.775 $Y=1.075 $X2=0 $Y2=0
cc_87 N_A_105_22#_c_75_n N_A1_c_230_n 0.0269594f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_88 N_A_105_22#_c_73_n N_A1_c_231_n 0.00184469f $X=1.775 $Y=1.075 $X2=0 $Y2=0
cc_89 N_A_105_22#_c_75_n N_A1_c_231_n 0.00147735f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_90 N_A_105_22#_c_73_n N_A1_c_232_n 0.00825902f $X=1.775 $Y=1.075 $X2=0 $Y2=0
cc_91 N_A_105_22#_c_74_n N_A1_c_232_n 9.48035e-19 $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_92 N_A_105_22#_c_75_n N_A1_c_232_n 0.00747875f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_93 N_A_105_22#_c_74_n N_A1_c_236_n 0.00731868f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_94 N_A_105_22#_c_74_n A1 0.104982f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_95 N_A_105_22#_c_75_n A1 0.025716f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_96 N_A_105_22#_c_74_n N_A0_M1005_g 0.00206802f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_97 N_A_105_22#_c_74_n N_A0_M1010_g 0.0139154f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_98 N_A_105_22#_c_75_n N_A0_M1010_g 0.0115019f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_99 N_A_105_22#_M1005_d A0 0.00489411f $X=1.8 $Y=2.17 $X2=0 $Y2=0
cc_100 N_A_105_22#_c_73_n A0 0.0124868f $X=1.775 $Y=1.075 $X2=0 $Y2=0
cc_101 N_A_105_22#_c_74_n A0 0.0818248f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_102 N_A_105_22#_c_75_n A0 0.00698325f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_103 N_A_105_22#_c_74_n N_A0_c_294_n 0.0155675f $X=2.185 $Y=2.375 $X2=0 $Y2=0
cc_104 N_A_105_22#_c_75_n N_A0_c_294_n 0.00611868f $X=1.94 $Y=0.87 $X2=0 $Y2=0
cc_105 N_A_105_22#_c_74_n N_A_488_106#_M1008_g 0.0012387f $X=2.185 $Y=2.375
+ $X2=0 $Y2=0
cc_106 N_A_105_22#_c_75_n N_A_488_106#_M1008_g 0.00172375f $X=1.94 $Y=0.87 $X2=0
+ $Y2=0
cc_107 N_A_105_22#_c_71_n N_X_c_389_n 0.0282825f $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_108 N_A_105_22#_c_117_p N_X_c_389_n 0.0105396f $X=0.9 $Y=1.075 $X2=0 $Y2=0
cc_109 N_A_105_22#_c_76_n N_X_c_389_n 0.0297165f $X=0.712 $Y=1.19 $X2=0 $Y2=0
cc_110 N_A_105_22#_M1006_g N_VPWR_c_402_n 0.0101853f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_105_22#_c_71_n N_VPWR_c_402_n 0.0108934f $X=0.735 $Y=1.355 $X2=0
+ $Y2=0
cc_112 N_A_105_22#_c_72_n N_VPWR_c_402_n 0.00139074f $X=0.735 $Y=1.355 $X2=0
+ $Y2=0
cc_113 N_A_105_22#_c_73_n N_VPWR_c_402_n 0.0038949f $X=1.775 $Y=1.075 $X2=0
+ $Y2=0
cc_114 N_A_105_22#_M1006_g N_VPWR_c_401_n 0.0129217f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_105_22#_M1006_g N_VPWR_c_408_n 0.00585385f $X=0.6 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_105_22#_c_73_n N_VGND_M1002_d 0.00642767f $X=1.775 $Y=1.075 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_105_22#_c_117_p N_VGND_M1002_d 0.00188388f $X=0.9 $Y=1.075 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_105_22#_c_72_n N_VGND_c_443_n 9.997e-19 $X=0.735 $Y=1.355 $X2=0 $Y2=0
cc_119 N_A_105_22#_c_73_n N_VGND_c_443_n 0.00639085f $X=1.775 $Y=1.075 $X2=0
+ $Y2=0
cc_120 N_A_105_22#_c_117_p N_VGND_c_443_n 0.0168254f $X=0.9 $Y=1.075 $X2=0 $Y2=0
cc_121 N_A_105_22#_c_76_n N_VGND_c_443_n 0.0128819f $X=0.712 $Y=1.19 $X2=0 $Y2=0
cc_122 N_A_105_22#_c_76_n N_VGND_c_447_n 0.009284f $X=0.712 $Y=1.19 $X2=0 $Y2=0
cc_123 N_A_105_22#_c_76_n N_VGND_c_448_n 0.0048178f $X=0.712 $Y=1.19 $X2=0 $Y2=0
cc_124 N_A_105_22#_c_73_n A_266_132# 0.00659274f $X=1.775 $Y=1.075 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_105_22#_c_75_n A_446_132# 7.79024e-19 $X=1.94 $Y=0.87 $X2=-0.19
+ $Y2=-0.245
cc_126 N_S_c_146_n N_A1_M1009_g 0.00444433f $X=2.905 $Y=2.97 $X2=0 $Y2=0
cc_127 N_S_c_148_n N_A1_M1009_g 3.706e-19 $X=2.99 $Y=2.13 $X2=0 $Y2=0
cc_128 N_S_c_149_n N_A1_M1009_g 0.00310312f $X=2.99 $Y=2.885 $X2=0 $Y2=0
cc_129 N_S_M1007_g N_A1_c_231_n 0.00133651f $X=1.255 $Y=0.87 $X2=0 $Y2=0
cc_130 N_S_M1007_g N_A1_c_232_n 0.0260657f $X=1.255 $Y=0.87 $X2=0 $Y2=0
cc_131 N_S_c_148_n N_A1_c_236_n 0.00190774f $X=2.99 $Y=2.13 $X2=0 $Y2=0
cc_132 N_S_c_146_n A1 0.0143563f $X=2.905 $Y=2.97 $X2=0 $Y2=0
cc_133 N_S_c_148_n A1 0.0346311f $X=2.99 $Y=2.13 $X2=0 $Y2=0
cc_134 N_S_c_149_n A1 0.0366856f $X=2.99 $Y=2.885 $X2=0 $Y2=0
cc_135 N_S_c_144_n N_A0_M1005_g 0.0341627f $X=1.275 $Y=2.01 $X2=0 $Y2=0
cc_136 N_S_c_138_n N_A0_M1005_g 7.80534e-19 $X=1.275 $Y=1.505 $X2=0 $Y2=0
cc_137 N_S_c_146_n N_A0_M1005_g 0.0042064f $X=2.905 $Y=2.97 $X2=0 $Y2=0
cc_138 N_S_c_139_n N_A0_M1010_g 0.00307675f $X=1.275 $Y=1.505 $X2=0 $Y2=0
cc_139 N_S_c_138_n A0 0.0823512f $X=1.275 $Y=1.505 $X2=0 $Y2=0
cc_140 N_S_c_139_n A0 0.00746485f $X=1.275 $Y=1.505 $X2=0 $Y2=0
cc_141 N_S_c_146_n A0 0.0146724f $X=2.905 $Y=2.97 $X2=0 $Y2=0
cc_142 N_S_c_137_n N_A0_c_294_n 0.0341627f $X=1.275 $Y=1.845 $X2=0 $Y2=0
cc_143 N_S_c_138_n N_A0_c_294_n 8.83096e-19 $X=1.275 $Y=1.505 $X2=0 $Y2=0
cc_144 N_S_c_148_n N_A_488_106#_c_332_n 0.00253186f $X=2.99 $Y=2.13 $X2=0 $Y2=0
cc_145 N_S_M1003_g N_A_488_106#_M1000_g 0.0292482f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_146 N_S_c_148_n N_A_488_106#_M1000_g 0.00701237f $X=2.99 $Y=2.13 $X2=0 $Y2=0
cc_147 N_S_c_149_n N_A_488_106#_M1000_g 0.0167846f $X=2.99 $Y=2.885 $X2=0 $Y2=0
cc_148 N_S_c_151_n N_A_488_106#_M1000_g 0.0115029f $X=3.685 $Y=1.845 $X2=0 $Y2=0
cc_149 N_S_M1003_g N_A_488_106#_c_335_n 0.016291f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_150 N_S_c_148_n N_A_488_106#_c_335_n 0.00758335f $X=2.99 $Y=2.13 $X2=0 $Y2=0
cc_151 N_S_c_151_n N_A_488_106#_c_335_n 0.0474594f $X=3.685 $Y=1.845 $X2=0 $Y2=0
cc_152 N_S_M1011_g N_A_488_106#_c_341_n 0.00358423f $X=3.595 $Y=2.38 $X2=0 $Y2=0
cc_153 N_S_c_150_n N_A_488_106#_c_341_n 8.63233e-19 $X=3.685 $Y=1.845 $X2=0
+ $Y2=0
cc_154 N_S_c_151_n N_A_488_106#_c_341_n 0.0143746f $X=3.685 $Y=1.845 $X2=0 $Y2=0
cc_155 N_S_M1003_g N_A_488_106#_c_336_n 0.0141992f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_156 N_S_M1003_g N_A_488_106#_c_337_n 0.00360909f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_157 N_S_M1011_g N_A_488_106#_c_337_n 0.00407587f $X=3.595 $Y=2.38 $X2=0 $Y2=0
cc_158 N_S_c_150_n N_A_488_106#_c_337_n 0.00353578f $X=3.685 $Y=1.845 $X2=0
+ $Y2=0
cc_159 N_S_c_151_n N_A_488_106#_c_337_n 0.031764f $X=3.685 $Y=1.845 $X2=0 $Y2=0
cc_160 N_S_M1003_g N_A_488_106#_c_338_n 0.00751856f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_161 N_S_c_150_n N_A_488_106#_c_338_n 0.00440081f $X=3.685 $Y=1.845 $X2=0
+ $Y2=0
cc_162 N_S_c_151_n N_A_488_106#_c_338_n 0.0158138f $X=3.685 $Y=1.845 $X2=0 $Y2=0
cc_163 N_S_M1003_g N_A_488_106#_c_339_n 0.0213806f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_164 N_S_c_151_n N_A_488_106#_c_339_n 0.00412429f $X=3.685 $Y=1.845 $X2=0
+ $Y2=0
cc_165 N_S_c_138_n N_VPWR_M1006_d 0.0039962f $X=1.275 $Y=1.505 $X2=-0.19
+ $Y2=-0.245
cc_166 N_S_M1004_g N_VPWR_c_402_n 0.00241231f $X=1.365 $Y=2.38 $X2=0 $Y2=0
cc_167 N_S_c_137_n N_VPWR_c_402_n 0.00190532f $X=1.275 $Y=1.845 $X2=0 $Y2=0
cc_168 N_S_c_138_n N_VPWR_c_402_n 0.0824087f $X=1.275 $Y=1.505 $X2=0 $Y2=0
cc_169 N_S_c_147_n N_VPWR_c_402_n 0.0149714f $X=1.36 $Y=2.97 $X2=0 $Y2=0
cc_170 N_S_M1011_g N_VPWR_c_403_n 0.00349123f $X=3.595 $Y=2.38 $X2=0 $Y2=0
cc_171 N_S_c_146_n N_VPWR_c_403_n 0.0146603f $X=2.905 $Y=2.97 $X2=0 $Y2=0
cc_172 N_S_c_149_n N_VPWR_c_403_n 0.0430535f $X=2.99 $Y=2.885 $X2=0 $Y2=0
cc_173 N_S_c_151_n N_VPWR_c_403_n 0.0195898f $X=3.685 $Y=1.845 $X2=0 $Y2=0
cc_174 N_S_M1004_g N_VPWR_c_404_n 2.80212e-19 $X=1.365 $Y=2.38 $X2=0 $Y2=0
cc_175 N_S_c_146_n N_VPWR_c_404_n 0.0992423f $X=2.905 $Y=2.97 $X2=0 $Y2=0
cc_176 N_S_c_147_n N_VPWR_c_404_n 0.0108172f $X=1.36 $Y=2.97 $X2=0 $Y2=0
cc_177 N_S_M1011_g N_VPWR_c_406_n 0.00347269f $X=3.595 $Y=2.38 $X2=0 $Y2=0
cc_178 N_S_M1011_g N_VPWR_c_401_n 0.00438782f $X=3.595 $Y=2.38 $X2=0 $Y2=0
cc_179 N_S_c_146_n N_VPWR_c_401_n 0.0639261f $X=2.905 $Y=2.97 $X2=0 $Y2=0
cc_180 N_S_c_147_n N_VPWR_c_401_n 0.00654547f $X=1.36 $Y=2.97 $X2=0 $Y2=0
cc_181 N_S_c_149_n A_518_434# 0.00371679f $X=2.99 $Y=2.885 $X2=-0.19 $Y2=-0.245
cc_182 N_S_M1007_g N_VGND_c_443_n 0.00713908f $X=1.255 $Y=0.87 $X2=0 $Y2=0
cc_183 N_S_M1003_g N_VGND_c_444_n 0.00635899f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_184 N_S_M1007_g N_VGND_c_445_n 0.00397346f $X=1.255 $Y=0.87 $X2=0 $Y2=0
cc_185 N_S_M1003_g N_VGND_c_446_n 0.00395058f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_186 N_S_M1007_g N_VGND_c_447_n 0.00459866f $X=1.255 $Y=0.87 $X2=0 $Y2=0
cc_187 N_S_M1003_g N_VGND_c_447_n 0.00459866f $X=3.595 $Y=0.87 $X2=0 $Y2=0
cc_188 N_A1_c_236_n N_A0_M1005_g 0.0105194f $X=2.605 $Y=1.845 $X2=0 $Y2=0
cc_189 A1 N_A0_M1005_g 3.00414e-19 $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_190 N_A1_c_230_n N_A0_M1010_g 0.00636498f $X=2.46 $Y=0.395 $X2=0 $Y2=0
cc_191 N_A1_c_231_n N_A0_M1010_g 0.00133993f $X=1.705 $Y=0.385 $X2=0 $Y2=0
cc_192 N_A1_c_232_n N_A0_M1010_g 0.0122971f $X=1.705 $Y=0.55 $X2=0 $Y2=0
cc_193 A1 N_A0_M1010_g 0.00434924f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_194 N_A1_M1009_g A0 0.00113765f $X=2.515 $Y=2.38 $X2=0 $Y2=0
cc_195 N_A1_c_232_n A0 0.00142189f $X=1.705 $Y=0.55 $X2=0 $Y2=0
cc_196 A1 A0 0.00121915f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_197 N_A1_c_232_n N_A0_c_294_n 0.00479482f $X=1.705 $Y=0.55 $X2=0 $Y2=0
cc_198 N_A1_c_236_n N_A0_c_294_n 0.0143801f $X=2.605 $Y=1.845 $X2=0 $Y2=0
cc_199 A1 N_A0_c_294_n 2.44928e-19 $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_200 N_A1_c_230_n N_A_488_106#_M1008_g 0.0012648f $X=2.46 $Y=0.395 $X2=0 $Y2=0
cc_201 N_A1_c_233_n N_A_488_106#_M1008_g 0.00271204f $X=2.597 $Y=0.535 $X2=0
+ $Y2=0
cc_202 A1 N_A_488_106#_M1008_g 0.0258986f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_203 A1 N_A_488_106#_c_332_n 0.00980408f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_204 N_A1_c_236_n N_A_488_106#_c_333_n 0.0138752f $X=2.605 $Y=1.845 $X2=0
+ $Y2=0
cc_205 A1 N_A_488_106#_c_333_n 0.00423024f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_206 N_A1_M1009_g N_A_488_106#_M1000_g 0.0201382f $X=2.515 $Y=2.38 $X2=0 $Y2=0
cc_207 N_A1_c_236_n N_A_488_106#_M1000_g 0.0205437f $X=2.605 $Y=1.845 $X2=0
+ $Y2=0
cc_208 A1 N_A_488_106#_M1000_g 0.00242105f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_209 A1 N_A_488_106#_c_335_n 0.0200078f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_210 A1 N_A_488_106#_c_339_n 0.0055947f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_211 A1 A_518_434# 0.00366783f $X=2.64 $Y=0.555 $X2=-0.19 $Y2=-0.245
cc_212 A1 N_VGND_M1008_d 0.00587549f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_213 N_A1_c_230_n N_VGND_c_443_n 0.00944439f $X=2.46 $Y=0.395 $X2=0 $Y2=0
cc_214 N_A1_c_231_n N_VGND_c_443_n 0.00224155f $X=1.705 $Y=0.385 $X2=0 $Y2=0
cc_215 N_A1_c_233_n N_VGND_c_444_n 0.0258431f $X=2.597 $Y=0.535 $X2=0 $Y2=0
cc_216 A1 N_VGND_c_444_n 0.0417382f $X=2.64 $Y=0.555 $X2=0 $Y2=0
cc_217 N_A1_c_230_n N_VGND_c_445_n 0.0603153f $X=2.46 $Y=0.395 $X2=0 $Y2=0
cc_218 N_A1_c_231_n N_VGND_c_445_n 0.00606749f $X=1.705 $Y=0.385 $X2=0 $Y2=0
cc_219 N_A1_c_233_n N_VGND_c_445_n 0.0197139f $X=2.597 $Y=0.535 $X2=0 $Y2=0
cc_220 N_A1_c_230_n N_VGND_c_447_n 0.0334616f $X=2.46 $Y=0.395 $X2=0 $Y2=0
cc_221 N_A1_c_231_n N_VGND_c_447_n 0.00851379f $X=1.705 $Y=0.385 $X2=0 $Y2=0
cc_222 N_A1_c_233_n N_VGND_c_447_n 0.0106914f $X=2.597 $Y=0.535 $X2=0 $Y2=0
cc_223 N_A0_M1010_g N_A_488_106#_M1008_g 0.0497281f $X=2.155 $Y=0.87 $X2=0 $Y2=0
cc_224 A0 A_288_434# 0.00431125f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_225 N_A0_M1010_g N_VGND_c_445_n 4.97633e-19 $X=2.155 $Y=0.87 $X2=0 $Y2=0
cc_226 N_A_488_106#_M1000_g N_VPWR_c_403_n 0.00318975f $X=3.055 $Y=2.38 $X2=0
+ $Y2=0
cc_227 N_A_488_106#_M1000_g N_VPWR_c_404_n 0.00160943f $X=3.055 $Y=2.38 $X2=0
+ $Y2=0
cc_228 N_A_488_106#_c_341_n N_VPWR_c_406_n 0.00770179f $X=4.03 $Y=2.435 $X2=0
+ $Y2=0
cc_229 N_A_488_106#_M1000_g N_VPWR_c_401_n 0.00162436f $X=3.055 $Y=2.38 $X2=0
+ $Y2=0
cc_230 N_A_488_106#_c_341_n N_VPWR_c_401_n 0.0148262f $X=4.03 $Y=2.435 $X2=0
+ $Y2=0
cc_231 N_A_488_106#_M1008_g N_VGND_c_444_n 0.002815f $X=2.515 $Y=0.87 $X2=0
+ $Y2=0
cc_232 N_A_488_106#_c_332_n N_VGND_c_444_n 0.011189f $X=2.98 $Y=1.295 $X2=0
+ $Y2=0
cc_233 N_A_488_106#_c_335_n N_VGND_c_444_n 0.0392168f $X=3.665 $Y=1.385 $X2=0
+ $Y2=0
cc_234 N_A_488_106#_M1008_g N_VGND_c_445_n 5.12641e-19 $X=2.515 $Y=0.87 $X2=0
+ $Y2=0
cc_235 N_A_488_106#_c_336_n N_VGND_c_446_n 0.00615429f $X=3.83 $Y=0.87 $X2=0
+ $Y2=0
cc_236 N_A_488_106#_c_336_n N_VGND_c_447_n 0.0113059f $X=3.83 $Y=0.87 $X2=0
+ $Y2=0
cc_237 N_X_c_389_n N_VPWR_c_402_n 0.0012507f $X=0.385 $Y=0.42 $X2=0 $Y2=0
cc_238 N_X_M1006_s N_VPWR_c_401_n 0.0040649f $X=0.26 $Y=1.835 $X2=0 $Y2=0
cc_239 N_X_c_389_n N_VPWR_c_401_n 0.0148849f $X=0.385 $Y=0.42 $X2=0 $Y2=0
cc_240 N_X_c_389_n N_VPWR_c_408_n 0.027134f $X=0.385 $Y=0.42 $X2=0 $Y2=0
cc_241 N_X_M1002_s N_VGND_c_447_n 0.00405061f $X=0.26 $Y=0.24 $X2=0 $Y2=0
cc_242 N_X_c_389_n N_VGND_c_447_n 0.0148849f $X=0.385 $Y=0.42 $X2=0 $Y2=0
cc_243 N_X_c_389_n N_VGND_c_448_n 0.027134f $X=0.385 $Y=0.42 $X2=0 $Y2=0
