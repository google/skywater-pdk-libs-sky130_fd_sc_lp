* File: sky130_fd_sc_lp__sdfbbn_2.spice
* Created: Wed Sep  2 10:33:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfbbn_2.pex.spice"
.subckt sky130_fd_sc_lp__sdfbbn_2  VNB VPB SCD D SCE CLK_N SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK_N	CLK_N
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1013 A_124_119# N_SCD_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1036 N_A_202_119#_M1036_d N_SCE_M1036_g A_124_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.09555 AS=0.0504 PD=0.875 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1019 A_323_119# N_D_M1019_g N_A_202_119#_M1036_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.09555 PD=0.84 PS=0.875 NRD=44.28 NRS=49.992 M=1 R=2.8
+ SA=75001.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_407_93#_M1004_g A_323_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.13335 AS=0.0882 PD=1.055 PS=0.84 NRD=47.136 NRS=44.28 M=1 R=2.8
+ SA=75001.8 SB=75001 A=0.063 P=1.14 MULT=1
MM1016 N_A_407_93#_M1016_d N_SCE_M1016_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.13335 PD=1.41 PS=1.055 NRD=0 NRS=54.276 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1049 N_A_840_95#_M1049_d N_CLK_N_M1049_g N_VGND_M1049_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.1533 PD=1.41 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75000.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_840_95#_M1010_g N_A_978_67#_M1010_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1218 AS=0.1449 PD=1.42 PS=1.53 NRD=5.712 NRS=17.136 M=1 R=2.8
+ SA=75000.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_1273_137#_M1011_d N_A_978_67#_M1011_g N_A_202_119#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1134 PD=0.7 PS=1.38 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1044 A_1359_137# N_A_840_95#_M1044_g N_A_1273_137#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.09765 AS=0.0588 PD=0.885 PS=0.7 NRD=50.712 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_1423_401#_M1017_g A_1359_137# VNB NSHORT L=0.15 W=0.42
+ AD=0.208158 AS=0.09765 PD=1.23226 PS=0.885 NRD=125.88 NRS=50.712 M=1 R=2.8
+ SA=75001.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1021 N_A_1670_93#_M1021_d N_SET_B_M1021_g N_VGND_M1017_d VNB NSHORT L=0.15
+ W=0.64 AD=0.096 AS=0.317192 PD=0.94 PS=1.87774 NRD=0 NRS=81.552 M=1 R=4.26667
+ SA=75001.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_1423_401#_M1029_d N_A_1273_137#_M1029_g N_A_1670_93#_M1021_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.14925 AS=0.096 PD=1.21 PS=0.94 NRD=33.408 NRS=0 M=1
+ R=4.26667 SA=75002.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1014 N_A_1670_93#_M1014_d N_A_1840_21#_M1014_g N_A_1423_401#_M1029_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1952 AS=0.14925 PD=1.89 PS=1.21 NRD=0 NRS=33.408 M=1
+ R=4.26667 SA=75002.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1046 A_2116_119# N_A_1423_401#_M1046_g N_VGND_M1046_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=23.436 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1022 N_A_2211_428#_M1022_d N_A_840_95#_M1022_g A_2116_119# VNB NSHORT L=0.15
+ W=0.64 AD=0.219955 AS=0.1152 PD=1.49132 PS=1 NRD=44.052 NRS=23.436 M=1
+ R=4.26667 SA=75000.7 SB=75002 A=0.096 P=1.58 MULT=1
MM1007 A_2367_163# N_A_978_67#_M1007_g N_A_2211_428#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.144345 PD=0.66 PS=0.978679 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_2415_137#_M1037_g A_2367_163# VNB NSHORT L=0.15 W=0.42
+ AD=0.143493 AS=0.0504 PD=1.10151 PS=0.66 NRD=81.9 NRS=18.564 M=1 R=2.8
+ SA=75001.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_2574_119#_M1030_d N_SET_B_M1030_g N_VGND_M1037_d VNB NSHORT L=0.15
+ W=0.64 AD=0.177775 AS=0.218657 PD=1.335 PS=1.67849 NRD=41.76 NRS=53.736 M=1
+ R=4.26667 SA=75001.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1047 N_A_2415_137#_M1047_d N_A_2211_428#_M1047_g N_A_2574_119#_M1030_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.125 AS=0.177775 PD=1.205 PS=1.335 NRD=8.436
+ NRS=41.76 M=1 R=4.26667 SA=75002.3 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1031 N_A_2574_119#_M1031_d N_A_1840_21#_M1031_g N_A_2415_137#_M1047_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1824 AS=0.125 PD=1.85 PS=1.205 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1032 N_VGND_M1032_d N_RESET_B_M1032_g N_A_1840_21#_M1032_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1032_d N_A_2415_137#_M1012_g N_Q_N_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1806 AS=0.1176 PD=1.6 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1041 N_VGND_M1041_d N_A_2415_137#_M1041_g N_Q_N_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2604 AS=0.1176 PD=2.3 PS=1.12 NRD=3.564 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1038 N_VGND_M1038_d N_A_2415_137#_M1038_g N_A_3289_47#_M1038_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_Q_M1003_d N_A_3289_47#_M1003_g N_VGND_M1038_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1806 PD=1.12 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1027 N_Q_M1003_d N_A_3289_47#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1048 N_VPWR_M1048_d N_SCD_M1048_g N_A_56_481#_M1048_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=24.6053 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1050 A_245_481# N_SCE_M1050_g N_VPWR_M1048_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1152 PD=0.88 PS=1 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1051 N_A_202_119#_M1051_d N_D_M1051_g A_245_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1344 AS=0.0768 PD=1.06 PS=0.88 NRD=18.4589 NRS=19.9955 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1015 N_A_56_481#_M1015_d N_A_407_93#_M1015_g N_A_202_119#_M1051_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=24.6053 M=1
+ R=4.26667 SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1028 N_A_407_93#_M1028_d N_SCE_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1728 AS=0.2846 PD=1.82 PS=3.18 NRD=0 NRS=119.934 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1025 N_A_840_95#_M1025_d N_CLK_N_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2784 AS=0.2368 PD=2.15 PS=2.02 NRD=52.3232 NRS=30.7714 M=1
+ R=4.26667 SA=75000.3 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_840_95#_M1008_g N_A_978_67#_M1008_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1728 AS=0.34125 PD=1.82 PS=2.96 NRD=0 NRS=147.179 M=1 R=4.26667
+ SA=75000.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1042 N_A_1273_137#_M1042_d N_A_840_95#_M1042_g N_A_202_119#_M1042_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0756 AS=0.1134 PD=0.78 PS=1.38 NRD=37.5088 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75006.3 A=0.063 P=1.14 MULT=1
MM1045 A_1375_463# N_A_978_67#_M1045_g N_A_1273_137#_M1042_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75005.8 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_1423_401#_M1018_g A_1375_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1792 AS=0.0504 PD=1.22333 PS=0.66 NRD=335.353 NRS=30.4759 M=1
+ R=2.8 SA=75001.1 SB=75005.4 A=0.063 P=1.14 MULT=1
MM1043 N_A_1423_401#_M1043_d N_SET_B_M1043_g N_VPWR_M1018_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1764 AS=0.3584 PD=1.26 PS=2.44667 NRD=32.8202 NRS=0 M=1 R=5.6
+ SA=75001.2 SB=75003.4 A=0.126 P=1.98 MULT=1
MM1033 A_1796_379# N_A_1273_137#_M1033_g N_A_1423_401#_M1043_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1008 AS=0.1764 PD=1.08 PS=1.26 NRD=15.2281 NRS=0 M=1 R=5.6
+ SA=75001.8 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_A_1840_21#_M1005_g A_1796_379# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.4452 AS=0.1008 PD=1.9 PS=1.08 NRD=38.6908 NRS=15.2281 M=1 R=5.6
+ SA=75002.2 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1039 A_2116_379# N_A_1423_401#_M1039_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.157937 AS=0.4452 PD=1.41 PS=1.9 NRD=31.1851 NRS=144.224 M=1 R=5.6
+ SA=75003.4 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1020 N_A_2211_428#_M1020_d N_A_978_67#_M1020_g A_2116_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1806 AS=0.157937 PD=1.6 PS=1.41 NRD=0 NRS=31.1851 M=1 R=5.6
+ SA=75003.1 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1009 A_2313_506# N_A_840_95#_M1009_g N_A_2211_428#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.14595 AS=0.0903 PD=1.115 PS=0.8 NRD=137.191 NRS=75.0373 M=1 R=2.8
+ SA=75003 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1035 N_VPWR_M1035_d N_A_2415_137#_M1035_g A_2313_506# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.119 AS=0.14595 PD=0.946667 PS=1.115 NRD=140.697 NRS=137.191 M=1
+ R=2.8 SA=75003.8 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1023 N_A_2415_137#_M1023_d N_SET_B_M1023_g N_VPWR_M1035_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.238 PD=1.12 PS=1.89333 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1000 A_2714_451# N_A_2211_428#_M1000_g N_A_2415_137#_M1023_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1008 AS=0.1176 PD=1.08 PS=1.12 NRD=15.2281 NRS=0 M=1 R=5.6
+ SA=75002.8 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1026 N_VPWR_M1026_d N_A_1840_21#_M1026_g A_2714_451# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2268 AS=0.1008 PD=2.22 PS=1.08 NRD=0 NRS=15.2281 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1040 N_VPWR_M1040_d N_RESET_B_M1040_g N_A_1840_21#_M1040_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.137128 AS=0.1728 PD=1.09137 PS=1.82 NRD=49.0136 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1040_d N_A_2415_137#_M1001_g N_Q_N_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.269972 AS=0.1764 PD=2.14863 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1024 N_VPWR_M1024_d N_A_2415_137#_M1024_g N_Q_N_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.378 AS=0.1764 PD=3.12 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4
+ SA=75000.9 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_2415_137#_M1006_g N_A_3289_47#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.137128 AS=0.1728 PD=1.09137 PS=1.82 NRD=25.3933 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_Q_M1002_d N_A_3289_47#_M1002_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.269972 PD=1.54 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1034 N_Q_M1002_d N_A_3289_47#_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX52_noxref VNB VPB NWDIODE A=35.0353 P=41.57
c_181 VNB 0 1.18451e-19 $X=0 $Y=0
c_349 VPB 0 1.58976e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfbbn_2.pxi.spice"
*
.ends
*
*
