* File: sky130_fd_sc_lp__sregsbp_1.spice
* Created: Fri Aug 28 11:33:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sregsbp_1.pex.spice"
.subckt sky130_fd_sc_lp__sregsbp_1  VNB VPB SCE D SCD CLK ASYNC VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* ASYNC	ASYNC
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1022 N_A_75_531#_M1022_d N_SCE_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 A_312_47# N_A_75_531#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1013 N_A_342_531#_M1013_d N_D_M1013_g A_312_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0504 PD=0.75 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1024 A_486_47# N_SCE_M1024_g N_A_342_531#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0693 PD=0.66 PS=0.75 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_SCD_M1025_g A_486_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1036 N_A_636_531#_M1036_d N_A_342_531#_M1036_g N_VGND_M1025_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_CLK_M1039_g N_A_761_357#_M1039_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1848 AS=0.2394 PD=1.28 PS=2.25 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1043 N_A_934_357#_M1043_d N_A_761_357#_M1043_g N_VGND_M1039_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.1848 PD=2.25 PS=1.28 NRD=0 NRS=11.424 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1032 N_A_1139_463#_M1032_d N_A_761_357#_M1032_g N_A_342_531#_M1032_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.09135 AS=0.1197 PD=0.855 PS=1.41 NRD=44.28 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1037 A_1319_119# N_A_934_357#_M1037_g N_A_1139_463#_M1032_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.09135 PD=0.63 PS=0.855 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1273_393#_M1001_g A_1319_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0914094 AS=0.0441 PD=0.824151 PS=0.63 NRD=34.284 NRS=14.28 M=1 R=2.8
+ SA=75001.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1038 A_1501_119# N_A_1139_463#_M1038_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.139291 PD=0.88 PS=1.25585 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_1273_393#_M1010_d N_ASYNC_M1010_g A_1501_119# VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 A_1825_125# N_A_1273_393#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.256 PD=0.88 PS=2.08 NRD=12.18 NRS=21.552 M=1 R=4.26667
+ SA=75000.3 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1027 N_A_1903_125#_M1027_d N_A_934_357#_M1027_g A_1825_125# VNB NSHORT L=0.15
+ W=0.64 AD=0.212226 AS=0.0768 PD=1.59396 PS=0.88 NRD=22.02 NRS=12.18 M=1
+ R=4.26667 SA=75000.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1021 A_2035_91# N_A_761_357#_M1021_g N_A_1903_125#_M1027_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.139274 PD=0.66 PS=1.04604 NRD=18.564 NRS=32.856 M=1
+ R=2.8 SA=75000.9 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_2083_65#_M1006_g A_2035_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.0905774 AS=0.0504 PD=0.820189 PS=0.66 NRD=34.284 NRS=18.564 M=1 R=2.8
+ SA=75001.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1040 A_2222_47# N_A_1903_125#_M1040_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.138023 PD=0.85 PS=1.24981 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_2083_65#_M1003_d N_ASYNC_M1003_g A_2222_47# VNB NSHORT L=0.15 W=0.64
+ AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75001.7
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 N_A_2456_451#_M1026_d N_A_2083_65#_M1026_g N_VGND_M1026_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_2083_65#_M1004_g N_Q_N_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1512 AS=0.2394 PD=1.2 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1016 N_Q_M1016_d N_A_2456_451#_M1016_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1512 PD=2.25 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1041 N_VPWR_M1041_d N_SCE_M1041_g N_A_75_531#_M1041_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=37.5088 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1000 A_264_531# N_SCE_M1000_g N_VPWR_M1041_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1020 N_A_342_531#_M1020_d N_D_M1020_g A_264_531# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1030 A_428_531# N_A_75_531#_M1030_g N_A_342_531#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0798 AS=0.0588 PD=0.8 PS=0.7 NRD=63.3158 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1028 N_VPWR_M1028_d N_SCD_M1028_g A_428_531# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0798 PD=0.78 PS=0.8 NRD=0 NRS=63.3158 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1031 N_A_636_531#_M1031_d N_A_342_531#_M1031_g N_VPWR_M1028_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=0 NRS=37.5088 M=1 R=2.8
+ SA=75002.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_CLK_M1005_g N_A_761_357#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_A_934_357#_M1029_d N_A_761_357#_M1029_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_A_1139_463#_M1009_d N_A_934_357#_M1009_g N_A_342_531#_M1009_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1017 A_1225_463# N_A_761_357#_M1017_g N_A_1139_463#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_VPWR_M1033_d N_A_1273_393#_M1033_g A_1225_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A_1139_463#_M1019_g N_A_1273_393#_M1019_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.255525 AS=0.2394 PD=1.635 PS=2.25 NRD=58.4302 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1034 N_A_1273_393#_M1034_d N_ASYNC_M1034_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2394 AS=0.255525 PD=2.25 PS=1.635 NRD=0 NRS=58.4302 M=1 R=5.6
+ SA=75000.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 A_1831_373# N_A_1273_393#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1638 AS=0.2394 PD=1.38 PS=2.25 NRD=32.8202 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1042 N_A_1903_125#_M1042_d N_A_761_357#_M1042_g A_1831_373# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1904 AS=0.1638 PD=1.64667 PS=1.38 NRD=0 NRS=32.8202 M=1 R=5.6
+ SA=75000.6 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1007 A_2042_451# N_A_934_357#_M1007_g N_A_1903_125#_M1042_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0952 PD=0.66 PS=0.823333 NRD=30.4759 NRS=56.2829 M=1
+ R=2.8 SA=75001.3 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_2083_65#_M1008_g A_2042_451# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0504 PD=0.876667 PS=0.66 NRD=105.533 NRS=30.4759 M=1 R=2.8
+ SA=75001.7 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1015 N_A_2083_65#_M1015_d N_A_1903_125#_M1015_g N_VPWR_M1008_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2352 PD=1.12 PS=1.75333 NRD=0 NRS=18.7544 M=1
+ R=5.6 SA=75001.3 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1035 N_VPWR_M1035_d N_ASYNC_M1035_g N_A_2083_65#_M1015_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.213973 AS=0.1176 PD=1.4927 PS=1.12 NRD=18.7544 NRS=0 M=1 R=5.6
+ SA=75001.7 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1023 N_A_2456_451#_M1023_d N_A_2083_65#_M1023_g N_VPWR_M1035_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.163027 PD=1.85 PS=1.1373 NRD=0 NRS=89.2607 M=1
+ R=4.26667 SA=75002.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_A_2083_65#_M1011_g N_Q_N_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.3591 PD=1.62 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1014 N_Q_M1014_d N_A_2456_451#_M1014_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.2268 PD=3.09 PS=1.62 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75000.7 SB=75000.2 A=0.189 P=2.82 MULT=1
DX44_noxref VNB VPB NWDIODE A=27.6402 P=33.39
c_155 VNB 0 4.80826e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__sregsbp_1.pxi.spice"
*
.ends
*
*
