* File: sky130_fd_sc_lp__nor4_m.spice
* Created: Fri Aug 28 10:57:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4_m.pex.spice"
.subckt sky130_fd_sc_lp__nor4_m  VNB VPB A B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1323 PD=0.7 PS=1.47 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.1092
+ AS=0.0588 PD=0.94 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.7 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_C_M1006_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1092 PD=0.7 PS=0.94 NRD=0 NRS=62.856 M=1 R=2.8 SA=75001.3 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_D_M1007_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1002 A_174_483# N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.1113 PD=0.66 PS=1.37 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1005 A_252_483# N_B_M1005_g A_174_483# VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=30.4759 NRS=30.4759 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_330_483# N_C_M1000_g A_252_483# VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=30.4759 NRS=30.4759 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_D_M1001_g A_330_483# VPB PHIGHVT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__nor4_m.pxi.spice"
*
.ends
*
*
