# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__dlrtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dlrtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.840000 1.015000 1.750000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.188600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.955000 0.255000 6.215000 0.585000 ;
        RECT 6.025000 0.585000 6.215000 1.085000 ;
        RECT 6.025000 1.085000 7.595000 1.255000 ;
        RECT 6.025000 1.765000 7.595000 1.935000 ;
        RECT 6.025000 1.935000 6.215000 3.075000 ;
        RECT 6.885000 0.255000 7.075000 1.085000 ;
        RECT 6.885000 1.935000 7.075000 3.075000 ;
        RECT 7.345000 1.255000 7.595000 1.765000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.210000 5.515000 2.130000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.920000 1.125000 2.150000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 7.680000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 7.870000 3.520000 ;
        RECT  1.375000 1.645000 2.215000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.095000  0.330000 0.625000 0.670000 ;
      RECT 0.095000  0.670000 0.365000 2.320000 ;
      RECT 0.095000  2.320000 1.125000 2.490000 ;
      RECT 0.095000  2.490000 0.365000 3.000000 ;
      RECT 0.535000  2.660000 0.785000 3.245000 ;
      RECT 0.795000  0.085000 1.125000 0.670000 ;
      RECT 0.955000  2.490000 1.125000 2.830000 ;
      RECT 0.955000  2.830000 2.010000 3.000000 ;
      RECT 1.295000  0.330000 1.495000 1.395000 ;
      RECT 1.295000  1.395000 1.920000 1.655000 ;
      RECT 1.295000  1.655000 1.505000 2.660000 ;
      RECT 1.675000  2.275000 2.835000 2.445000 ;
      RECT 1.675000  2.445000 2.010000 2.830000 ;
      RECT 1.745000  1.825000 2.270000 2.105000 ;
      RECT 1.900000  0.735000 2.110000 1.055000 ;
      RECT 1.900000  1.055000 3.375000 1.225000 ;
      RECT 2.100000  1.225000 2.270000 1.825000 ;
      RECT 2.290000  0.085000 2.620000 0.875000 ;
      RECT 2.325000  2.615000 2.655000 3.245000 ;
      RECT 2.505000  1.405000 2.835000 2.275000 ;
      RECT 2.820000  0.255000 3.735000 0.495000 ;
      RECT 2.820000  0.495000 2.990000 1.055000 ;
      RECT 3.045000  1.225000 3.375000 2.075000 ;
      RECT 3.170000  0.665000 3.725000 0.885000 ;
      RECT 3.190000  2.245000 3.725000 2.885000 ;
      RECT 3.545000  0.885000 3.725000 1.065000 ;
      RECT 3.545000  1.065000 4.775000 1.235000 ;
      RECT 3.545000  1.235000 3.725000 2.245000 ;
      RECT 3.950000  1.405000 4.280000 2.300000 ;
      RECT 3.950000  2.300000 5.855000 2.470000 ;
      RECT 4.070000  0.085000 4.400000 0.895000 ;
      RECT 4.525000  1.235000 4.775000 1.515000 ;
      RECT 4.590000  0.255000 4.920000 0.725000 ;
      RECT 4.590000  0.725000 5.115000 0.870000 ;
      RECT 4.590000  0.870000 5.855000 0.895000 ;
      RECT 4.590000  2.640000 4.920000 3.245000 ;
      RECT 4.945000  0.895000 5.855000 1.040000 ;
      RECT 5.090000  2.470000 5.310000 3.075000 ;
      RECT 5.445000  0.085000 5.775000 0.700000 ;
      RECT 5.480000  2.640000 5.810000 3.245000 ;
      RECT 5.685000  1.040000 5.855000 1.425000 ;
      RECT 5.685000  1.425000 7.175000 1.595000 ;
      RECT 5.685000  1.595000 5.855000 2.300000 ;
      RECT 6.385000  0.085000 6.715000 0.915000 ;
      RECT 6.385000  2.105000 6.715000 3.245000 ;
      RECT 7.245000  0.085000 7.575000 0.915000 ;
      RECT 7.245000  2.105000 7.575000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrtn_4
END LIBRARY
