* File: sky130_fd_sc_lp__xnor2_0.spice
* Created: Wed Sep  2 10:39:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor2_0.pex.spice"
.subckt sky130_fd_sc_lp__xnor2_0  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 A_110_177# N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_143_487#_M1001_d N_B_M1001_g A_110_177# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_300_60#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_300_60#_M1009_d N_B_M1009_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_143_487#_M1002_g N_A_300_60#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_143_487#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_143_487#_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1984 AS=0.0896 PD=1.26 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1005 A_383_487# N_A_M1005_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1984 PD=0.85 PS=1.26 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75001.4 SB=75001
+ A=0.096 P=1.58 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g A_383_487# VPB PHIGHVT L=0.15 W=0.64 AD=0.096
+ AS=0.0672 PD=0.94 PS=0.85 NRD=6.1464 NRS=15.3857 M=1 R=4.26667 SA=75001.8
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_143_487#_M1008_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.096 PD=1.81 PS=0.94 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__xnor2_0.pxi.spice"
*
.ends
*
*
