* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
X0 Q a_857_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_857_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_599_47# a_414_47# a_671_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_671_47# a_857_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_49_70# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 Q a_857_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND a_857_21# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_828_469# a_857_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 Q a_857_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_651_469# a_267_464# a_671_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_671_47# a_267_464# a_779_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_779_47# a_857_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_414_47# a_267_464# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 Q a_857_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR a_857_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND a_49_70# a_599_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_414_47# a_267_464# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_671_47# a_414_47# a_828_469# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 VPWR a_857_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_857_21# a_671_47# a_1083_73# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR a_49_70# a_651_469# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VGND GATE a_267_464# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1083_73# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 VGND a_857_21# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VPWR GATE a_267_464# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_49_70# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
