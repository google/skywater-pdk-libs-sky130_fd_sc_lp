# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrbp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrbp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.500000 1.180000 0.835000 1.850000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.160000 1.715000 7.615000 2.890000 ;
        RECT 7.445000 0.265000 7.820000 0.685000 ;
        RECT 7.445000 0.685000 7.615000 1.715000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.370000 1.850000 9.960000 2.890000 ;
        RECT 9.630000 0.350000 9.960000 0.810000 ;
        RECT 9.725000 0.810000 9.960000 1.850000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.795000 1.920000 8.125000 2.890000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.675000 1.850000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.540000  0.445000 1.000000 ;
      RECT 0.115000  1.000000  0.285000 2.075000 ;
      RECT 0.115000  2.075000  0.605000 2.515000 ;
      RECT 0.115000  2.515000  2.155000 2.685000 ;
      RECT 0.115000  2.685000  0.605000 3.065000 ;
      RECT 0.805000  2.865000  1.135000 3.245000 ;
      RECT 0.905000  0.085000  1.235000 1.000000 ;
      RECT 1.335000  2.075000  1.665000 2.165000 ;
      RECT 1.335000  2.165000  2.975000 2.335000 ;
      RECT 1.695000  0.540000  2.025000 1.000000 ;
      RECT 1.825000  2.685000  2.155000 3.065000 ;
      RECT 1.855000  1.000000  2.025000 2.165000 ;
      RECT 2.255000  0.265000  2.585000 0.785000 ;
      RECT 2.255000  0.785000  4.040000 0.955000 ;
      RECT 2.255000  0.955000  2.425000 1.655000 ;
      RECT 2.255000  1.655000  2.625000 1.985000 ;
      RECT 2.645000  1.135000  2.975000 1.345000 ;
      RECT 2.645000  1.345000  4.000000 1.465000 ;
      RECT 2.805000  1.465000  4.000000 1.675000 ;
      RECT 2.805000  1.675000  2.975000 2.165000 ;
      RECT 2.905000  2.515000  3.235000 3.245000 ;
      RECT 3.045000  0.085000  3.375000 0.605000 ;
      RECT 3.670000  1.675000  4.000000 2.895000 ;
      RECT 3.670000  2.895000  4.900000 3.065000 ;
      RECT 3.710000  0.775000  4.040000 0.785000 ;
      RECT 3.710000  0.955000  4.040000 1.105000 ;
      RECT 4.180000  1.815000  4.510000 2.715000 ;
      RECT 4.220000  0.265000  4.550000 0.515000 ;
      RECT 4.220000  0.515000  5.250000 0.685000 ;
      RECT 4.220000  0.685000  4.390000 1.815000 ;
      RECT 4.570000  0.865000  4.900000 1.195000 ;
      RECT 4.730000  1.195000  4.900000 2.895000 ;
      RECT 5.080000  0.685000  5.250000 0.865000 ;
      RECT 5.080000  0.865000  6.040000 1.035000 ;
      RECT 5.140000  1.345000  5.470000 1.715000 ;
      RECT 5.140000  1.715000  6.390000 1.885000 ;
      RECT 5.365000  2.065000  5.695000 3.245000 ;
      RECT 5.430000  0.085000  5.680000 0.685000 ;
      RECT 5.710000  1.035000  6.040000 1.535000 ;
      RECT 5.910000  0.305000  6.390000 0.685000 ;
      RECT 6.015000  1.885000  6.390000 2.855000 ;
      RECT 6.220000  0.685000  6.390000 1.365000 ;
      RECT 6.220000  1.365000  7.265000 1.535000 ;
      RECT 6.220000  1.535000  6.390000 1.715000 ;
      RECT 6.625000  1.715000  6.955000 3.245000 ;
      RECT 6.700000  0.085000  7.030000 0.685000 ;
      RECT 6.935000  0.865000  7.265000 1.365000 ;
      RECT 8.050000  0.350000  8.380000 0.990000 ;
      RECT 8.050000  0.990000  9.475000 1.160000 ;
      RECT 8.310000  1.160000  8.640000 2.890000 ;
      RECT 8.840000  0.085000  9.170000 0.810000 ;
      RECT 8.840000  1.850000  9.170000 3.245000 ;
      RECT 9.145000  1.160000  9.475000 1.660000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrbp_lp
END LIBRARY
