* File: sky130_fd_sc_lp__o311a_lp.pex.spice
* Created: Wed Sep  2 10:23:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311A_LP%A_84_115# 1 2 3 10 12 15 19 22 24 27 28 31
+ 32 33 36 38 45 46 48 50
r92 45 50 3.95216 $w=2.32e-07 $l=1.12161e-07 $layer=LI1_cond $X=3.665 $Y=2.1
+ $X2=3.602 $Y2=2.185
r93 44 45 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.665 $Y=1.07
+ $X2=3.665 $Y2=2.1
r94 38 44 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.58 $Y=0.905
+ $X2=3.665 $Y2=1.07
r95 38 40 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.58 $Y=0.905
+ $X2=3.315 $Y2=0.905
r96 37 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=2.185
+ $X2=2.46 $Y2=2.185
r97 36 50 2.49072 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.455 $Y=2.185
+ $X2=3.602 $Y2=2.185
r98 36 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.455 $Y=2.185
+ $X2=2.625 $Y2=2.185
r99 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=2.185
+ $X2=2.46 $Y2=2.185
r100 32 33 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=2.295 $Y=2.185
+ $X2=0.81 $Y2=2.185
r101 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.725 $Y=2.1
+ $X2=0.81 $Y2=2.185
r102 31 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=2.1
+ $X2=0.725 $Y2=1.935
r103 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=1.43 $X2=0.615 $Y2=1.43
r104 25 46 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.63 $Y=1.755
+ $X2=0.63 $Y2=1.935
r105 25 27 10.404 $w=3.58e-07 $l=3.25e-07 $layer=LI1_cond $X=0.63 $Y=1.755
+ $X2=0.63 $Y2=1.43
r106 23 28 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=0.6 $Y=1.755
+ $X2=0.6 $Y2=1.43
r107 23 24 33.13 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.6 $Y=1.755 $X2=0.6
+ $Y2=1.935
r108 22 28 12.8232 $w=3.6e-07 $l=8e-08 $layer=POLY_cond $X=0.6 $Y=1.35 $X2=0.6
+ $Y2=1.43
r109 15 24 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.56 $Y=2.595
+ $X2=0.56 $Y2=1.935
r110 10 22 25.8164 $w=3.6e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=1.2
+ $X2=0.675 $Y2=1.35
r111 10 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=1.2
+ $X2=0.855 $Y2=0.915
r112 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.2
+ $X2=0.495 $Y2=0.915
r113 3 50 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=3.4
+ $Y=2.095 $X2=3.54 $Y2=2.265
r114 2 48 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=2.095 $X2=2.46 $Y2=2.265
r115 1 40 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.705 $X2=3.315 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%A1 3 9 10 11 12 15 17
c41 12 0 4.22402e-20 $X=1.2 $Y=1.665
r42 15 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.755
+ $X2=1.155 $Y2=1.92
r43 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.755
+ $X2=1.155 $Y2=1.59
r44 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.755 $X2=1.155 $Y2=1.755
r45 12 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.155 $Y=1.665
+ $X2=1.155 $Y2=1.755
r46 11 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.245 $Y=1.35
+ $X2=1.245 $Y2=1.59
r47 10 11 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=1.267 $Y=1.2
+ $X2=1.267 $Y2=1.35
r48 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.29 $Y=0.915 $X2=1.29
+ $Y2=1.2
r49 3 18 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.165 $Y=2.595
+ $X2=1.165 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%A2 3 7 9 12
c38 7 0 1.60424e-19 $X=1.72 $Y=0.915
r39 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.755
+ $X2=1.695 $Y2=1.92
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.755
+ $X2=1.695 $Y2=1.59
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.695
+ $Y=1.755 $X2=1.695 $Y2=1.755
r42 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.755
r43 7 14 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.72 $Y=0.915
+ $X2=1.72 $Y2=1.59
r44 3 15 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.655 $Y=2.595
+ $X2=1.655 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%A3 3 7 9 12
c37 9 0 1.54746e-19 $X=2.16 $Y=1.665
r38 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.715
+ $X2=2.235 $Y2=1.88
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.715
+ $X2=2.235 $Y2=1.55
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.715 $X2=2.235 $Y2=1.715
r41 7 14 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.31 $Y=0.915
+ $X2=2.31 $Y2=1.55
r42 3 15 177.644 $w=2.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.195 $Y=2.595
+ $X2=2.195 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%B1 3 7 9 12 13
c37 13 0 1.06774e-19 $X=2.775 $Y=1.755
c38 7 0 1.66705e-19 $X=2.74 $Y=0.915
r39 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.755
+ $X2=2.775 $Y2=1.92
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.755
+ $X2=2.775 $Y2=1.59
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.775
+ $Y=1.755 $X2=2.775 $Y2=1.755
r42 9 13 4.20486 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.64 $Y=1.735
+ $X2=2.775 $Y2=1.735
r43 7 14 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.74 $Y=0.915
+ $X2=2.74 $Y2=1.59
r44 3 15 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.735 $Y=2.595
+ $X2=2.735 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%C1 1 3 8 12 14 17 18 19
c36 19 0 1.98852e-19 $X=3.315 $Y=1.59
c37 18 0 1.30142e-19 $X=3.315 $Y=1.755
r38 17 20 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.755
+ $X2=3.315 $Y2=1.92
r39 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.755
+ $X2=3.315 $Y2=1.59
r40 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.315
+ $Y=1.755 $X2=3.315 $Y2=1.755
r41 14 18 6.07369 $w=3.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.12 $Y=1.735
+ $X2=3.315 $Y2=1.735
r42 10 12 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.1 $Y=1.275
+ $X2=3.225 $Y2=1.275
r43 8 20 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.275 $Y=2.595
+ $X2=3.275 $Y2=1.92
r44 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.225 $Y=1.35
+ $X2=3.225 $Y2=1.275
r45 4 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.225 $Y=1.35
+ $X2=3.225 $Y2=1.59
r46 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=1.2 $X2=3.1
+ $Y2=1.275
r47 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.1 $Y=1.2 $X2=3.1
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%X 1 2 12 13 14 15 26
r22 19 26 0.40085 $w=3.43e-07 $l=1.2e-08 $layer=LI1_cond $X=0.272 $Y=0.913
+ $X2=0.272 $Y2=0.925
r23 15 28 7.10983 $w=3.43e-07 $l=1.24e-07 $layer=LI1_cond $X=0.272 $Y=0.961
+ $X2=0.272 $Y2=1.085
r24 15 26 1.20255 $w=3.43e-07 $l=3.6e-08 $layer=LI1_cond $X=0.272 $Y=0.961
+ $X2=0.272 $Y2=0.925
r25 15 19 1.23595 $w=3.43e-07 $l=3.7e-08 $layer=LI1_cond $X=0.272 $Y=0.876
+ $X2=0.272 $Y2=0.913
r26 14 15 10.7227 $w=3.43e-07 $l=3.21e-07 $layer=LI1_cond $X=0.272 $Y=0.555
+ $X2=0.272 $Y2=0.876
r27 13 28 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.185 $Y=2.115
+ $X2=0.185 $Y2=1.085
r28 12 13 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.28
+ $X2=0.28 $Y2=2.115
r29 2 12 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.095 $X2=0.295 $Y2=2.28
r30 1 15 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.705 $X2=0.28 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%VPWR 1 2 11 15 18 19 20 30 31 34
r45 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.825 $Y2=3.33
r53 22 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 18 27 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33 $X2=3
+ $Y2=3.33
r58 17 30 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33 $X2=3
+ $Y2=3.33
r60 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=3.33
r61 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.78
r62 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=3.33
r63 9 11 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=2.78
r64 2 15 600 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=2.095 $X2=3 $Y2=2.78
r65 1 11 600 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.095 $X2=0.825 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%VGND 1 2 9 13 16 17 18 24 30 31 34
r39 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 31 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r42 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.015
+ $Y2=0
r43 28 30 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=2.18 $Y=0 $X2=3.6
+ $Y2=0
r44 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.015
+ $Y2=0
r46 24 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r47 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r48 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r50 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r51 16 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r52 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.03
+ $Y2=0
r53 15 26 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.68
+ $Y2=0
r54 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.03
+ $Y2=0
r55 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0
r56 11 13 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0.85
r57 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=0.085
+ $X2=1.03 $Y2=0
r58 7 9 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=1.03 $Y=0.085 $X2=1.03
+ $Y2=0.885
r59 2 13 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.795
+ $Y=0.705 $X2=2.015 $Y2=0.85
r60 1 9 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.93 $Y=0.705
+ $X2=1.07 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_LP%A_273_141# 1 2 7 11 14
c33 7 0 9.20776e-20 $X=2.36 $Y=1.285
r34 14 15 16.296 $w=2.77e-07 $l=3.7e-07 $layer=LI1_cond $X=1.505 $Y=0.915
+ $X2=1.505 $Y2=1.285
r35 9 11 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.525 $Y=1.2
+ $X2=2.525 $Y2=0.915
r36 8 15 3.59349 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=1.285
+ $X2=1.505 $Y2=1.285
r37 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.36 $Y=1.285
+ $X2=2.525 $Y2=1.2
r38 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.36 $Y=1.285 $X2=1.67
+ $Y2=1.285
r39 2 11 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.705 $X2=2.525 $Y2=0.915
r40 1 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.705 $X2=1.505 $Y2=0.915
.ends

