* File: sky130_fd_sc_lp__ebufn_lp.pex.spice
* Created: Fri Aug 28 10:32:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EBUFN_LP%A 3 7 11 15 17 18 22 23
r38 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.655
+ $Y=1.41 $X2=0.655 $Y2=1.41
r39 17 18 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.662 $Y=1.665
+ $X2=0.662 $Y2=2.035
r40 17 23 8.51806 $w=3.43e-07 $l=2.55e-07 $layer=LI1_cond $X=0.662 $Y=1.665
+ $X2=0.662 $Y2=1.41
r41 13 22 92.2311 $w=2.7e-07 $l=5.94559e-07 $layer=POLY_cond $X=0.895 $Y=1.915
+ $X2=0.7 $Y2=1.41
r42 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.895 $Y=1.915
+ $X2=0.895 $Y2=2.735
r43 9 22 31.5348 $w=2.7e-07 $l=2.64953e-07 $layer=POLY_cond $X=0.895 $Y=1.245
+ $X2=0.7 $Y2=1.41
r44 9 11 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.895 $Y=1.245
+ $X2=0.895 $Y2=0.865
r45 5 22 31.5348 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.41
+ $X2=0.7 $Y2=1.41
r46 5 7 194.851 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.535 $Y=1.41
+ $X2=0.535 $Y2=0.865
r47 1 22 92.2311 $w=2.7e-07 $l=5.94559e-07 $layer=POLY_cond $X=0.505 $Y=1.915
+ $X2=0.7 $Y2=1.41
r48 1 3 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.505 $Y=1.915
+ $X2=0.505 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP%A_242_237# 1 2 9 10 13 16 17 18 20 21 22 25
+ 29 33 34 36
c75 29 0 1.11563e-19 $X=4.04 $Y=2.15
c76 13 0 1.26037e-19 $X=1.375 $Y=1.35
r77 31 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.12 $Y=1.005
+ $X2=4.04 $Y2=0.92
r78 31 34 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.12 $Y=1.005
+ $X2=4.12 $Y2=1.985
r79 29 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=2.15
+ $X2=4.04 $Y2=1.985
r80 23 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.835
+ $X2=4.04 $Y2=0.92
r81 23 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.04 $Y=0.835
+ $X2=4.04 $Y2=0.465
r82 21 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=0.92
+ $X2=4.04 $Y2=0.92
r83 21 22 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.875 $Y=0.92
+ $X2=2.915 $Y2=0.92
r84 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.83 $Y=0.835
+ $X2=2.915 $Y2=0.92
r85 19 20 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.83 $Y=0.425
+ $X2=2.83 $Y2=0.835
r86 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.745 $Y=0.34
+ $X2=2.83 $Y2=0.425
r87 17 18 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.745 $Y=0.34
+ $X2=1.735 $Y2=0.34
r88 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.65 $Y=0.425
+ $X2=1.735 $Y2=0.34
r89 15 16 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.65 $Y=0.425
+ $X2=1.65 $Y2=1.185
r90 13 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.35
+ $X2=1.375 $Y2=1.185
r91 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.375
+ $Y=1.35 $X2=1.375 $Y2=1.35
r92 10 16 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.35
+ $X2=1.65 $Y2=1.185
r93 10 12 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.565 $Y=1.35
+ $X2=1.375 $Y2=1.35
r94 9 36 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.465 $Y=0.655
+ $X2=1.465 $Y2=1.185
r95 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.9
+ $Y=2.005 $X2=4.04 $Y2=2.15
r96 1 25 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.04 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP%A_29_483# 1 2 9 11 15 18 21 24 25 26 29 33
+ 37 41
c69 29 0 1.26037e-19 $X=2.07 $Y=1.51
r70 33 35 10.2717 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.305 $Y=0.855
+ $X2=0.305 $Y2=1.075
r71 30 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.51
+ $X2=2.235 $Y2=1.51
r72 30 38 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.07 $Y=1.51
+ $X2=1.855 $Y2=1.51
r73 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.51 $X2=2.07 $Y2=1.51
r74 27 29 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.07 $Y=1.685
+ $X2=2.07 $Y2=1.51
r75 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.905 $Y=1.77
+ $X2=2.07 $Y2=1.685
r76 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.905 $Y=1.77
+ $X2=1.175 $Y2=1.77
r77 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=1.855
+ $X2=1.175 $Y2=1.77
r78 23 24 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.09 $Y=1.855
+ $X2=1.09 $Y2=2.395
r79 22 37 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=2.48
+ $X2=0.29 $Y2=2.48
r80 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.005 $Y=2.48
+ $X2=1.09 $Y2=2.395
r81 21 22 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.005 $Y=2.48
+ $X2=0.455 $Y2=2.48
r82 18 37 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.21 $Y=2.395
+ $X2=0.29 $Y2=2.48
r83 18 35 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=0.21 $Y=2.395
+ $X2=0.21 $Y2=1.075
r84 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.5 $Y=1.675 $X2=2.5
+ $Y2=2.465
r85 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.425 $Y=1.6
+ $X2=2.5 $Y2=1.675
r86 11 41 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.425 $Y=1.6
+ $X2=2.235 $Y2=1.6
r87 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=1.51
r88 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=0.655
r89 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=2.415 $X2=0.29 $Y2=2.56
r90 1 33 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.655 $X2=0.32 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP%TE_B 3 5 6 9 13 15 17 19 21 23 26 28 29
c56 15 0 1.11563e-19 $X=3.825 $Y=1.175
r57 33 35 27.8843 $w=2.42e-07 $l=1.4e-07 $layer=POLY_cond $X=3.465 $Y=1.34
+ $X2=3.605 $Y2=1.34
r58 32 33 5.97521 $w=2.42e-07 $l=3e-08 $layer=POLY_cond $X=3.435 $Y=1.34
+ $X2=3.465 $Y2=1.34
r59 28 29 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.605 $Y=1.295
+ $X2=3.605 $Y2=1.665
r60 28 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.605
+ $Y=1.34 $X2=3.605 $Y2=1.34
r61 24 26 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.825 $Y=1.82
+ $X2=4.085 $Y2=1.82
r62 23 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.085 $Y=1.745
+ $X2=4.085 $Y2=1.82
r63 22 23 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.085 $Y=1.325
+ $X2=4.085 $Y2=1.745
r64 19 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.825 $Y=1.895
+ $X2=3.825 $Y2=1.82
r65 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.825 $Y=1.895
+ $X2=3.825 $Y2=2.325
r66 15 22 51.7851 $w=2.42e-07 $l=3.26497e-07 $layer=POLY_cond $X=3.825 $Y=1.175
+ $X2=4.085 $Y2=1.325
r67 15 35 43.8182 $w=2.42e-07 $l=2.91033e-07 $layer=POLY_cond $X=3.825 $Y=1.175
+ $X2=3.605 $Y2=1.34
r68 15 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.825 $Y=1.175
+ $X2=3.825 $Y2=0.445
r69 11 33 13.9682 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.465 $Y=1.175
+ $X2=3.465 $Y2=1.34
r70 11 13 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.465 $Y=1.175
+ $X2=3.465 $Y2=0.445
r71 7 32 13.9682 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.435 $Y=1.505
+ $X2=3.435 $Y2=1.34
r72 7 9 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.435 $Y=1.505
+ $X2=3.435 $Y2=2.325
r73 5 32 21.8618 $w=2.42e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.36 $Y=1.25
+ $X2=3.435 $Y2=1.34
r74 5 6 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.36 $Y=1.25
+ $X2=2.965 $Y2=1.25
r75 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.89 $Y=1.325
+ $X2=2.965 $Y2=1.25
r76 1 3 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.89 $Y=1.325
+ $X2=2.89 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP%VPWR 1 2 9 13 20 21 22 31 40 41 44
r42 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 41 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 38 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.27 $Y=3.33
+ $X2=3.105 $Y2=3.33
r46 38 40 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.27 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 37 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r50 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.94 $Y=3.33
+ $X2=3.105 $Y2=3.33
r52 31 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.94 $Y=3.33 $X2=2.64
+ $Y2=3.33
r53 30 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 26 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 25 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 22 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 20 29 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.51 $Y2=3.33
r62 19 33 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=1.51 $Y2=3.33
r64 16 18 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.105 $Y=2.465
+ $X2=3.105 $Y2=2.95
r65 13 16 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.105 $Y=1.98
+ $X2=3.105 $Y2=2.465
r66 11 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=3.245
+ $X2=3.105 $Y2=3.33
r67 11 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.105 $Y=3.245
+ $X2=3.105 $Y2=2.95
r68 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=3.245 $X2=1.51
+ $Y2=3.33
r69 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.51 $Y=3.245
+ $X2=1.51 $Y2=2.56
r70 2 18 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.835 $X2=3.105 $Y2=2.95
r71 2 16 600 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.835 $X2=3.105 $Y2=2.465
r72 2 13 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.835 $X2=3.105 $Y2=1.98
r73 1 9 300 $w=1.7e-07 $l=6.08194e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=2.415 $X2=1.51 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP%Z 1 2 7 8 9 10 11 31
r31 20 31 2.12386 $w=5.81e-07 $l=1.47916e-07 $layer=LI1_cond $X=2.58 $Y=2.025
+ $X2=2.437 $Y2=2.035
r32 19 26 13.9195 $w=4.47e-07 $l=6.72964e-07 $layer=LI1_cond $X=2.58 $Y=1.35
+ $X2=2.07 $Y2=0.972
r33 11 40 2.83477 $w=5.81e-07 $l=1.35e-07 $layer=LI1_cond $X=2.437 $Y=2.775
+ $X2=2.437 $Y2=2.91
r34 10 11 7.76936 $w=5.81e-07 $l=3.7e-07 $layer=LI1_cond $X=2.437 $Y=2.405
+ $X2=2.437 $Y2=2.775
r35 10 34 4.51463 $w=5.81e-07 $l=2.15e-07 $layer=LI1_cond $X=2.437 $Y=2.405
+ $X2=2.437 $Y2=2.19
r36 9 34 2.4778 $w=5.81e-07 $l=1.18e-07 $layer=LI1_cond $X=2.437 $Y=2.072
+ $X2=2.437 $Y2=2.19
r37 9 31 0.776936 $w=5.81e-07 $l=3.7e-08 $layer=LI1_cond $X=2.437 $Y=2.072
+ $X2=2.437 $Y2=2.035
r38 9 20 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=2.58 $Y=1.987
+ $X2=2.58 $Y2=2.025
r39 8 9 10.6025 $w=3.48e-07 $l=3.22e-07 $layer=LI1_cond $X=2.58 $Y=1.665
+ $X2=2.58 $Y2=1.987
r40 7 19 1.63758 $w=4.47e-07 $l=9.53939e-08 $layer=LI1_cond $X=2.64 $Y=1.28
+ $X2=2.58 $Y2=1.35
r41 7 8 9.87808 $w=3.48e-07 $l=3e-07 $layer=LI1_cond $X=2.58 $Y=1.365 $X2=2.58
+ $Y2=1.665
r42 7 19 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=2.58 $Y=1.365
+ $X2=2.58 $Y2=1.35
r43 2 40 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.835 $X2=2.285 $Y2=2.91
r44 2 34 400 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.835 $X2=2.285 $Y2=2.19
r45 1 26 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.235 $X2=2.07 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_LP%VGND 1 2 9 15 17 19 24 31 32 35 38
r47 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r50 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r51 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.25
+ $Y2=0
r52 29 31 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=4.08
+ $Y2=0
r53 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.23
+ $Y2=0
r56 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.68
+ $Y2=0
r57 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.25
+ $Y2=0
r58 24 27 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=3.085 $Y=0
+ $X2=1.68 $Y2=0
r59 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r60 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.23
+ $Y2=0
r62 19 21 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r63 17 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r64 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r65 13 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r66 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0.44
r67 9 11 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.23 $Y=0.38 $X2=1.23
+ $Y2=0.85
r68 7 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085 $X2=1.23
+ $Y2=0
r69 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.38
r70 2 15 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.25 $Y2=0.44
r71 1 11 182 $w=1.7e-07 $l=3.43948e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.655 $X2=1.23 $Y2=0.85
r72 1 9 182 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.655 $X2=1.23 $Y2=0.38
.ends

