# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__iso1n_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__iso1n_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.189000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.910000 1.395000 2.580000 1.750000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.160000 1.160000 1.990000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.445200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 0.465000 3.755000 3.075000 ;
    END
  END X
  PIN KAGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.070000 0.440000 3.770000 0.670000 ;
    END
  END KAGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.120000  0.430000 0.365000 0.885000 ;
      RECT 0.125000  0.885000 0.370000 2.160000 ;
      RECT 0.125000  2.160000 1.700000 2.330000 ;
      RECT 0.345000  2.330000 0.590000 2.820000 ;
      RECT 0.885000  0.430000 1.515000 0.885000 ;
      RECT 1.190000  2.500000 1.520000 3.245000 ;
      RECT 1.370000  1.315000 1.700000 2.160000 ;
      RECT 1.735000  0.430000 2.065000 0.885000 ;
      RECT 1.870000  0.885000 2.065000 1.055000 ;
      RECT 1.870000  1.055000 3.225000 1.225000 ;
      RECT 2.095000  1.955000 3.225000 2.125000 ;
      RECT 2.095000  2.125000 2.305000 2.880000 ;
      RECT 2.525000  0.430000 3.155000 0.885000 ;
      RECT 2.525000  2.295000 2.910000 3.245000 ;
      RECT 2.895000  1.225000 3.225000 1.955000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 0.935000  0.470000 1.105000 0.640000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.295000  0.470000 1.465000 0.640000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 2.575000  0.470000 2.745000 0.640000 ;
      RECT 2.935000  0.470000 3.105000 0.640000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__iso1n_lp
END LIBRARY
