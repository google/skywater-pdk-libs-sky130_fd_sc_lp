* File: sky130_fd_sc_lp__clkinv_16.pex.spice
* Created: Wed Sep  2 09:40:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINV_16%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55
+ 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131 135 139 143
+ 147 151 155 159 161 220 223 231 236 241 246 251 256 261 266 270
r374 267 270 0.692933 $w=2.3e-07 $l=1.08e-06 $layer=MET1_cond $X=9.3 $Y=1.295
+ $X2=10.38 $Y2=1.295
r375 266 270 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.38 $Y=1.295
+ $X2=10.38 $Y2=1.295
r376 266 267 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.3 $Y=1.295
+ $X2=9.3 $Y2=1.295
r377 262 267 0.708973 $w=2.3e-07 $l=1.105e-06 $layer=MET1_cond $X=8.195 $Y=1.295
+ $X2=9.3 $Y2=1.295
r378 261 262 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.195 $Y=1.295
+ $X2=8.195 $Y2=1.295
r379 257 262 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.335 $Y=1.295
+ $X2=8.195 $Y2=1.295
r380 256 257 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.335 $Y=1.295
+ $X2=7.335 $Y2=1.295
r381 252 257 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.475 $Y=1.295
+ $X2=7.335 $Y2=1.295
r382 251 252 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.475 $Y=1.295
+ $X2=6.475 $Y2=1.295
r383 241 242 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.755 $Y=1.295
+ $X2=4.755 $Y2=1.295
r384 237 242 0.554988 $w=2.3e-07 $l=8.65e-07 $layer=MET1_cond $X=3.89 $Y=1.295
+ $X2=4.755 $Y2=1.295
r385 236 237 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.89 $Y=1.295
+ $X2=3.89 $Y2=1.295
r386 232 237 0.548572 $w=2.3e-07 $l=8.55e-07 $layer=MET1_cond $X=3.035 $Y=1.295
+ $X2=3.89 $Y2=1.295
r387 231 232 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.035 $Y=1.295
+ $X2=3.035 $Y2=1.295
r388 227 232 0.702557 $w=2.3e-07 $l=1.095e-06 $layer=MET1_cond $X=1.94 $Y=1.295
+ $X2=3.035 $Y2=1.295
r389 224 227 0.692933 $w=2.3e-07 $l=1.08e-06 $layer=MET1_cond $X=0.86 $Y=1.295
+ $X2=1.94 $Y2=1.295
r390 223 227 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.94 $Y=1.295
+ $X2=1.94 $Y2=1.295
r391 223 224 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.86 $Y=1.295
+ $X2=0.86 $Y2=1.295
r392 218 220 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=10.38 $Y=1.46
+ $X2=10.555 $Y2=1.46
r393 216 218 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=10.125 $Y=1.46
+ $X2=10.38 $Y2=1.46
r394 215 216 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=9.695 $Y=1.46
+ $X2=10.125 $Y2=1.46
r395 214 215 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=9.265 $Y=1.46
+ $X2=9.695 $Y2=1.46
r396 213 266 1.23877 $w=1.623e-06 $l=1.65e-07 $layer=LI1_cond $X=9.732 $Y=1.46
+ $X2=9.732 $Y2=1.295
r397 213 218 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=10.38
+ $Y=1.46 $X2=10.38 $Y2=1.46
r398 212 214 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=9.02 $Y=1.46
+ $X2=9.265 $Y2=1.46
r399 212 213 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.02
+ $Y=1.46 $X2=9.02 $Y2=1.46
r400 210 212 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=8.835 $Y=1.46
+ $X2=9.02 $Y2=1.46
r401 209 210 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.405 $Y=1.46
+ $X2=8.835 $Y2=1.46
r402 207 209 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.195 $Y=1.46
+ $X2=8.405 $Y2=1.46
r403 207 261 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.195
+ $Y=1.46 $X2=8.195 $Y2=1.46
r404 205 207 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=7.975 $Y=1.46
+ $X2=8.195 $Y2=1.46
r405 204 205 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.545 $Y=1.46
+ $X2=7.975 $Y2=1.46
r406 202 204 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.335 $Y=1.46
+ $X2=7.545 $Y2=1.46
r407 202 256 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.335
+ $Y=1.46 $X2=7.335 $Y2=1.46
r408 200 202 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=7.115 $Y=1.46
+ $X2=7.335 $Y2=1.46
r409 199 200 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.685 $Y=1.46
+ $X2=7.115 $Y2=1.46
r410 197 199 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.475 $Y=1.46
+ $X2=6.685 $Y2=1.46
r411 197 251 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.475
+ $Y=1.46 $X2=6.475 $Y2=1.46
r412 195 197 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=6.255 $Y=1.46
+ $X2=6.475 $Y2=1.46
r413 194 195 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.825 $Y=1.46
+ $X2=6.255 $Y2=1.46
r414 192 194 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.61 $Y=1.46
+ $X2=5.825 $Y2=1.46
r415 192 246 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.61
+ $Y=1.46 $X2=5.61 $Y2=1.46
r416 190 192 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.395 $Y=1.46
+ $X2=5.61 $Y2=1.46
r417 189 190 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.965 $Y=1.46
+ $X2=5.395 $Y2=1.46
r418 187 189 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.755 $Y=1.46
+ $X2=4.965 $Y2=1.46
r419 187 241 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.46 $X2=4.755 $Y2=1.46
r420 185 187 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=4.535 $Y=1.46
+ $X2=4.755 $Y2=1.46
r421 184 185 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.105 $Y=1.46
+ $X2=4.535 $Y2=1.46
r422 182 184 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.89 $Y=1.46
+ $X2=4.105 $Y2=1.46
r423 182 236 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.46 $X2=3.89 $Y2=1.46
r424 180 182 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.675 $Y=1.46
+ $X2=3.89 $Y2=1.46
r425 179 180 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.245 $Y=1.46
+ $X2=3.675 $Y2=1.46
r426 177 179 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.035 $Y=1.46
+ $X2=3.245 $Y2=1.46
r427 177 231 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.035
+ $Y=1.46 $X2=3.035 $Y2=1.46
r428 175 177 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.815 $Y=1.46
+ $X2=3.035 $Y2=1.46
r429 174 175 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.385 $Y=1.46
+ $X2=2.815 $Y2=1.46
r430 172 174 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=1.46
+ $X2=2.385 $Y2=1.46
r431 170 172 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.955 $Y=1.46
+ $X2=2.22 $Y2=1.46
r432 169 170 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.525 $Y=1.46
+ $X2=1.955 $Y2=1.46
r433 168 169 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.095 $Y=1.46
+ $X2=1.525 $Y2=1.46
r434 167 223 1.17376 $w=1.713e-06 $l=1.65e-07 $layer=LI1_cond $X=1.447 $Y=1.46
+ $X2=1.447 $Y2=1.295
r435 167 172 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.22
+ $Y=1.46 $X2=2.22 $Y2=1.46
r436 166 168 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.86 $Y=1.46
+ $X2=1.095 $Y2=1.46
r437 166 167 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.86
+ $Y=1.46 $X2=0.86 $Y2=1.46
r438 163 166 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.665 $Y=1.46
+ $X2=0.86 $Y2=1.46
r439 161 252 0.554988 $w=2.3e-07 $l=8.65e-07 $layer=MET1_cond $X=5.61 $Y=1.295
+ $X2=6.475 $Y2=1.295
r440 161 242 0.548572 $w=2.3e-07 $l=8.55e-07 $layer=MET1_cond $X=5.61 $Y=1.295
+ $X2=4.755 $Y2=1.295
r441 161 246 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.295
r442 157 220 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.555 $Y=1.625
+ $X2=10.555 $Y2=1.46
r443 157 159 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=10.555 $Y=1.625
+ $X2=10.555 $Y2=2.465
r444 153 216 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.125 $Y=1.625
+ $X2=10.125 $Y2=1.46
r445 153 155 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=10.125 $Y=1.625
+ $X2=10.125 $Y2=2.465
r446 149 215 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.695 $Y=1.625
+ $X2=9.695 $Y2=1.46
r447 149 151 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.695 $Y=1.625
+ $X2=9.695 $Y2=2.465
r448 145 214 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.265 $Y=1.625
+ $X2=9.265 $Y2=1.46
r449 145 147 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.265 $Y=1.625
+ $X2=9.265 $Y2=2.465
r450 141 210 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.835 $Y=1.625
+ $X2=8.835 $Y2=1.46
r451 141 143 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.835 $Y=1.625
+ $X2=8.835 $Y2=2.465
r452 137 210 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.835 $Y=1.295
+ $X2=8.835 $Y2=1.46
r453 137 139 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=8.835 $Y=1.295
+ $X2=8.835 $Y2=0.56
r454 133 209 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.405 $Y=1.625
+ $X2=8.405 $Y2=1.46
r455 133 135 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.405 $Y=1.625
+ $X2=8.405 $Y2=2.465
r456 129 209 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.405 $Y=1.295
+ $X2=8.405 $Y2=1.46
r457 129 131 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=8.405 $Y=1.295
+ $X2=8.405 $Y2=0.56
r458 125 205 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.975 $Y=1.625
+ $X2=7.975 $Y2=1.46
r459 125 127 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.975 $Y=1.625
+ $X2=7.975 $Y2=2.465
r460 121 205 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.975 $Y=1.295
+ $X2=7.975 $Y2=1.46
r461 121 123 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=7.975 $Y=1.295
+ $X2=7.975 $Y2=0.56
r462 117 204 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.545 $Y=1.625
+ $X2=7.545 $Y2=1.46
r463 117 119 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.545 $Y=1.625
+ $X2=7.545 $Y2=2.465
r464 113 204 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.545 $Y=1.295
+ $X2=7.545 $Y2=1.46
r465 113 115 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=7.545 $Y=1.295
+ $X2=7.545 $Y2=0.56
r466 109 200 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.115 $Y=1.625
+ $X2=7.115 $Y2=1.46
r467 109 111 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.115 $Y=1.625
+ $X2=7.115 $Y2=2.465
r468 105 200 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.115 $Y=1.295
+ $X2=7.115 $Y2=1.46
r469 105 107 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=7.115 $Y=1.295
+ $X2=7.115 $Y2=0.56
r470 101 199 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.685 $Y=1.625
+ $X2=6.685 $Y2=1.46
r471 101 103 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.685 $Y=1.625
+ $X2=6.685 $Y2=2.465
r472 97 199 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.685 $Y=1.295
+ $X2=6.685 $Y2=1.46
r473 97 99 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=6.685 $Y=1.295
+ $X2=6.685 $Y2=0.56
r474 93 195 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.625
+ $X2=6.255 $Y2=1.46
r475 93 95 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.255 $Y=1.625
+ $X2=6.255 $Y2=2.465
r476 89 195 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.295
+ $X2=6.255 $Y2=1.46
r477 89 91 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=6.255 $Y=1.295
+ $X2=6.255 $Y2=0.56
r478 85 194 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.625
+ $X2=5.825 $Y2=1.46
r479 85 87 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.825 $Y=1.625
+ $X2=5.825 $Y2=2.465
r480 81 194 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.295
+ $X2=5.825 $Y2=1.46
r481 81 83 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=5.825 $Y=1.295
+ $X2=5.825 $Y2=0.56
r482 77 190 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.625
+ $X2=5.395 $Y2=1.46
r483 77 79 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.395 $Y=1.625
+ $X2=5.395 $Y2=2.465
r484 73 190 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.295
+ $X2=5.395 $Y2=1.46
r485 73 75 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=5.395 $Y=1.295
+ $X2=5.395 $Y2=0.56
r486 69 189 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.625
+ $X2=4.965 $Y2=1.46
r487 69 71 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.965 $Y=1.625
+ $X2=4.965 $Y2=2.465
r488 65 189 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.295
+ $X2=4.965 $Y2=1.46
r489 65 67 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=4.965 $Y=1.295
+ $X2=4.965 $Y2=0.56
r490 61 185 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.535 $Y=1.625
+ $X2=4.535 $Y2=1.46
r491 61 63 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.535 $Y=1.625
+ $X2=4.535 $Y2=2.465
r492 57 185 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.535 $Y=1.295
+ $X2=4.535 $Y2=1.46
r493 57 59 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=4.535 $Y=1.295
+ $X2=4.535 $Y2=0.56
r494 53 184 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=1.46
r495 53 55 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=2.465
r496 49 184 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.295
+ $X2=4.105 $Y2=1.46
r497 49 51 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=4.105 $Y=1.295
+ $X2=4.105 $Y2=0.56
r498 45 180 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.675 $Y=1.625
+ $X2=3.675 $Y2=1.46
r499 45 47 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.675 $Y=1.625
+ $X2=3.675 $Y2=2.465
r500 41 180 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.675 $Y=1.295
+ $X2=3.675 $Y2=1.46
r501 41 43 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=3.675 $Y=1.295
+ $X2=3.675 $Y2=0.56
r502 37 179 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.245 $Y=1.625
+ $X2=3.245 $Y2=1.46
r503 37 39 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.245 $Y=1.625
+ $X2=3.245 $Y2=2.465
r504 33 179 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.245 $Y=1.295
+ $X2=3.245 $Y2=1.46
r505 33 35 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=3.245 $Y=1.295
+ $X2=3.245 $Y2=0.56
r506 29 175 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.625
+ $X2=2.815 $Y2=1.46
r507 29 31 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.815 $Y=1.625
+ $X2=2.815 $Y2=2.465
r508 25 175 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.295
+ $X2=2.815 $Y2=1.46
r509 25 27 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=2.815 $Y=1.295
+ $X2=2.815 $Y2=0.56
r510 21 174 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.625
+ $X2=2.385 $Y2=1.46
r511 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.385 $Y=1.625
+ $X2=2.385 $Y2=2.465
r512 17 174 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.295
+ $X2=2.385 $Y2=1.46
r513 17 19 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=2.385 $Y=1.295
+ $X2=2.385 $Y2=0.56
r514 13 170 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.625
+ $X2=1.955 $Y2=1.46
r515 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.955 $Y=1.625
+ $X2=1.955 $Y2=2.465
r516 9 169 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.625
+ $X2=1.525 $Y2=1.46
r517 9 11 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.525 $Y=1.625
+ $X2=1.525 $Y2=2.465
r518 5 168 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.625
+ $X2=1.095 $Y2=1.46
r519 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.095 $Y=1.625
+ $X2=1.095 $Y2=2.465
r520 1 163 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.625
+ $X2=0.665 $Y2=1.46
r521 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.665 $Y=1.625
+ $X2=0.665 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 42 46
+ 50 56 62 68 74 78 82 88 94 100 106 110 114 118 120 124 125 127 128 130 131 132
+ 133 135 136 138 139 140 141 142 148 163 178 184 187 190 193 196 200
r228 199 200 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r229 196 197 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r230 193 194 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r231 187 188 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r232 184 185 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r233 182 200 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r234 182 197 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r235 181 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r236 179 196 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.04 $Y=3.33
+ $X2=9.91 $Y2=3.33
r237 179 181 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.04 $Y=3.33
+ $X2=10.32 $Y2=3.33
r238 178 199 4.00962 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.64 $Y=3.33
+ $X2=10.84 $Y2=3.33
r239 178 181 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.64 $Y=3.33
+ $X2=10.32 $Y2=3.33
r240 177 197 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r241 176 177 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r242 174 177 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r243 173 174 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r244 171 174 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r245 171 194 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r246 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r247 168 193 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.47 $Y2=3.33
r248 168 170 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r249 167 194 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r250 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r251 164 190 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.74 $Y=3.33
+ $X2=5.61 $Y2=3.33
r252 164 166 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.74 $Y=3.33
+ $X2=6 $Y2=3.33
r253 163 193 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.34 $Y=3.33
+ $X2=6.47 $Y2=3.33
r254 163 166 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.34 $Y=3.33
+ $X2=6 $Y2=3.33
r255 161 162 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r256 159 162 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r257 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r258 156 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r259 156 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r260 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r261 153 187 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.17 $Y2=3.33
r262 153 155 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.64 $Y2=3.33
r263 152 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r264 152 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r265 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r266 149 184 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.44 $Y=3.33
+ $X2=1.31 $Y2=3.33
r267 149 151 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r268 148 187 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=2.17 $Y2=3.33
r269 148 151 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r270 146 185 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r271 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r272 142 167 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r273 142 162 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r274 142 190 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r275 140 176 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=8.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r276 140 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.92 $Y=3.33
+ $X2=9.05 $Y2=3.33
r277 138 173 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=7.92 $Y2=3.33
r278 138 139 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=8.19 $Y2=3.33
r279 137 176 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.32 $Y=3.33
+ $X2=8.88 $Y2=3.33
r280 137 139 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.32 $Y=3.33
+ $X2=8.19 $Y2=3.33
r281 135 170 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r282 135 136 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.2 $Y=3.33
+ $X2=7.33 $Y2=3.33
r283 134 173 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.46 $Y=3.33
+ $X2=7.92 $Y2=3.33
r284 134 136 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.46 $Y=3.33
+ $X2=7.33 $Y2=3.33
r285 132 161 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.62 $Y=3.33
+ $X2=4.56 $Y2=3.33
r286 132 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.62 $Y=3.33
+ $X2=4.75 $Y2=3.33
r287 130 158 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.6 $Y2=3.33
r288 130 131 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.89 $Y2=3.33
r289 129 161 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=4.56 $Y2=3.33
r290 129 131 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=3.89 $Y2=3.33
r291 127 155 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=2.64 $Y2=3.33
r292 127 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=3.03 $Y2=3.33
r293 126 158 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r294 126 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=3.03 $Y2=3.33
r295 124 145 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.32 $Y=3.33
+ $X2=0.24 $Y2=3.33
r296 124 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.32 $Y=3.33
+ $X2=0.45 $Y2=3.33
r297 120 123 38.4148 $w=2.53e-07 $l=8.5e-07 $layer=LI1_cond $X=10.767 $Y=2.04
+ $X2=10.767 $Y2=2.89
r298 118 199 3.1676 $w=2.55e-07 $l=1.15888e-07 $layer=LI1_cond $X=10.767
+ $Y=3.245 $X2=10.84 $Y2=3.33
r299 118 123 16.0438 $w=2.53e-07 $l=3.55e-07 $layer=LI1_cond $X=10.767 $Y=3.245
+ $X2=10.767 $Y2=2.89
r300 114 117 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=9.91 $Y=2.04
+ $X2=9.91 $Y2=2.89
r301 112 196 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.91 $Y=3.245
+ $X2=9.91 $Y2=3.33
r302 112 117 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=9.91 $Y=3.245
+ $X2=9.91 $Y2=2.89
r303 111 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.18 $Y=3.33
+ $X2=9.05 $Y2=3.33
r304 110 196 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.78 $Y=3.33
+ $X2=9.91 $Y2=3.33
r305 110 111 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=9.78 $Y=3.33
+ $X2=9.18 $Y2=3.33
r306 106 109 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=9.05 $Y=2.04
+ $X2=9.05 $Y2=2.89
r307 104 141 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.05 $Y=3.245
+ $X2=9.05 $Y2=3.33
r308 104 109 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=9.05 $Y=3.245
+ $X2=9.05 $Y2=2.89
r309 100 103 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=8.19 $Y=2.04
+ $X2=8.19 $Y2=2.89
r310 98 139 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.19 $Y=3.245
+ $X2=8.19 $Y2=3.33
r311 98 103 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=8.19 $Y=3.245
+ $X2=8.19 $Y2=2.89
r312 94 97 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=7.33 $Y=2.04
+ $X2=7.33 $Y2=2.89
r313 92 136 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=3.245
+ $X2=7.33 $Y2=3.33
r314 92 97 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=7.33 $Y=3.245
+ $X2=7.33 $Y2=2.89
r315 88 91 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=6.47 $Y=2.04
+ $X2=6.47 $Y2=2.89
r316 86 193 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=3.33
r317 86 91 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=2.89
r318 82 85 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=5.61 $Y=2.04
+ $X2=5.61 $Y2=2.89
r319 80 190 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.61 $Y=3.245
+ $X2=5.61 $Y2=3.33
r320 80 85 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=5.61 $Y=3.245
+ $X2=5.61 $Y2=2.89
r321 79 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=4.75 $Y2=3.33
r322 78 190 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=5.61 $Y2=3.33
r323 78 79 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.48 $Y=3.33 $X2=4.88
+ $Y2=3.33
r324 74 77 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=4.75 $Y=2.04
+ $X2=4.75 $Y2=2.89
r325 72 133 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=3.33
r326 72 77 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=2.89
r327 68 71 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=3.89 $Y=2.04
+ $X2=3.89 $Y2=2.89
r328 66 131 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=3.245
+ $X2=3.89 $Y2=3.33
r329 66 71 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=3.89 $Y=3.245
+ $X2=3.89 $Y2=2.89
r330 62 65 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=3.03 $Y=2.04
+ $X2=3.03 $Y2=2.89
r331 60 128 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=3.33
r332 60 65 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=2.89
r333 56 59 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=2.17 $Y=2.04
+ $X2=2.17 $Y2=2.89
r334 54 187 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r335 54 59 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.89
r336 50 53 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=1.31 $Y=2.04
+ $X2=1.31 $Y2=2.89
r337 48 184 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=3.245
+ $X2=1.31 $Y2=3.33
r338 48 53 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=1.31 $Y=3.245
+ $X2=1.31 $Y2=2.89
r339 47 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.45 $Y2=3.33
r340 46 184 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.18 $Y=3.33
+ $X2=1.31 $Y2=3.33
r341 46 47 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.18 $Y=3.33 $X2=0.58
+ $Y2=3.33
r342 42 45 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=0.45 $Y=2.04
+ $X2=0.45 $Y2=2.89
r343 40 125 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.45 $Y=3.245
+ $X2=0.45 $Y2=3.33
r344 40 45 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=0.45 $Y=3.245
+ $X2=0.45 $Y2=2.89
r345 13 123 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.835 $X2=10.77 $Y2=2.89
r346 13 120 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.835 $X2=10.77 $Y2=2.04
r347 12 117 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=9.77
+ $Y=1.835 $X2=9.91 $Y2=2.89
r348 12 114 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=9.77
+ $Y=1.835 $X2=9.91 $Y2=2.04
r349 11 109 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=8.91
+ $Y=1.835 $X2=9.05 $Y2=2.89
r350 11 106 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=8.91
+ $Y=1.835 $X2=9.05 $Y2=2.04
r351 10 103 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=8.05
+ $Y=1.835 $X2=8.19 $Y2=2.89
r352 10 100 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=8.05
+ $Y=1.835 $X2=8.19 $Y2=2.04
r353 9 97 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=7.19
+ $Y=1.835 $X2=7.33 $Y2=2.89
r354 9 94 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.19
+ $Y=1.835 $X2=7.33 $Y2=2.04
r355 8 91 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=6.33
+ $Y=1.835 $X2=6.47 $Y2=2.89
r356 8 88 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=6.33
+ $Y=1.835 $X2=6.47 $Y2=2.04
r357 7 85 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=5.47
+ $Y=1.835 $X2=5.61 $Y2=2.89
r358 7 82 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.47
+ $Y=1.835 $X2=5.61 $Y2=2.04
r359 6 77 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=4.61
+ $Y=1.835 $X2=4.75 $Y2=2.89
r360 6 74 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=4.61
+ $Y=1.835 $X2=4.75 $Y2=2.04
r361 5 71 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.75
+ $Y=1.835 $X2=3.89 $Y2=2.89
r362 5 68 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.75
+ $Y=1.835 $X2=3.89 $Y2=2.04
r363 4 65 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=1.835 $X2=3.03 $Y2=2.89
r364 4 62 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=1.835 $X2=3.03 $Y2=2.04
r365 3 59 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.835 $X2=2.17 $Y2=2.89
r366 3 56 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.835 $X2=2.17 $Y2=2.04
r367 2 53 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=1.17
+ $Y=1.835 $X2=1.31 $Y2=2.89
r368 2 50 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.17
+ $Y=1.835 $X2=1.31 $Y2=2.04
r369 1 45 400 $w=1.7e-07 $l=1.12517e-06 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.835 $X2=0.45 $Y2=2.89
r370 1 42 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.835 $X2=0.45 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 63 65 67 70 78 86 96 106 116 123 133 143 153 163 171 172
r237 171 176 37.8976 $w=2.58e-07 $l=8.55e-07 $layer=LI1_cond $X=10.34 $Y=2.035
+ $X2=10.34 $Y2=2.89
r238 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.34 $Y=2.035
+ $X2=10.34 $Y2=2.035
r239 164 172 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=9.48 $Y=2.035
+ $X2=10.34 $Y2=2.035
r240 163 168 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=9.482 $Y=2.035
+ $X2=9.482 $Y2=2.89
r241 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.48 $Y=2.035
+ $X2=9.48 $Y2=2.035
r242 157 164 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=8.62 $Y=2.035
+ $X2=9.48 $Y2=2.035
r243 156 160 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=8.622 $Y=2.035
+ $X2=8.622 $Y2=2.89
r244 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.62 $Y=2.035
+ $X2=8.62 $Y2=2.035
r245 153 156 66.6609 $w=2.53e-07 $l=1.475e-06 $layer=LI1_cond $X=8.622 $Y=0.56
+ $X2=8.622 $Y2=2.035
r246 147 157 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=7.76 $Y=2.035
+ $X2=8.62 $Y2=2.035
r247 146 150 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=7.762 $Y=2.035
+ $X2=7.762 $Y2=2.89
r248 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.76 $Y=2.035
+ $X2=7.76 $Y2=2.035
r249 143 146 66.6609 $w=2.53e-07 $l=1.475e-06 $layer=LI1_cond $X=7.762 $Y=0.56
+ $X2=7.762 $Y2=2.035
r250 137 147 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.9 $Y=2.035
+ $X2=7.76 $Y2=2.035
r251 136 140 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=6.902 $Y=2.035
+ $X2=6.902 $Y2=2.89
r252 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.9 $Y=2.035
+ $X2=6.9 $Y2=2.035
r253 133 136 66.6609 $w=2.53e-07 $l=1.475e-06 $layer=LI1_cond $X=6.902 $Y=0.56
+ $X2=6.902 $Y2=2.035
r254 127 137 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=6.04 $Y=2.035
+ $X2=6.9 $Y2=2.035
r255 126 130 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=6.042 $Y=2.035
+ $X2=6.042 $Y2=2.89
r256 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.04 $Y=2.035
+ $X2=6.04 $Y2=2.035
r257 123 126 66.6609 $w=2.53e-07 $l=1.475e-06 $layer=LI1_cond $X=6.042 $Y=0.56
+ $X2=6.042 $Y2=2.035
r258 116 120 37.8976 $w=2.58e-07 $l=8.55e-07 $layer=LI1_cond $X=5.18 $Y=2.035
+ $X2=5.18 $Y2=2.89
r259 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.18 $Y=2.035
+ $X2=5.18 $Y2=2.035
r260 110 117 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=4.32 $Y=2.035
+ $X2=5.18 $Y2=2.035
r261 109 113 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=4.322 $Y=2.035
+ $X2=4.322 $Y2=2.89
r262 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.32 $Y=2.035
+ $X2=4.32 $Y2=2.035
r263 106 109 66.6609 $w=2.53e-07 $l=1.475e-06 $layer=LI1_cond $X=4.322 $Y=0.56
+ $X2=4.322 $Y2=2.035
r264 100 110 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=3.46 $Y=2.035
+ $X2=4.32 $Y2=2.035
r265 99 103 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=3.462 $Y=2.035
+ $X2=3.462 $Y2=2.89
r266 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.46 $Y=2.035
+ $X2=3.46 $Y2=2.035
r267 96 99 66.6609 $w=2.53e-07 $l=1.475e-06 $layer=LI1_cond $X=3.462 $Y=0.56
+ $X2=3.462 $Y2=2.035
r268 90 100 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=2.6 $Y=2.035
+ $X2=3.46 $Y2=2.035
r269 89 93 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=2.602 $Y=2.035
+ $X2=2.602 $Y2=2.89
r270 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.6 $Y=2.035
+ $X2=2.6 $Y2=2.035
r271 86 89 66.6609 $w=2.53e-07 $l=1.475e-06 $layer=LI1_cond $X=2.602 $Y=0.56
+ $X2=2.602 $Y2=2.035
r272 79 90 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=1.74 $Y=2.035
+ $X2=2.6 $Y2=2.035
r273 78 83 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=1.742 $Y=2.035
+ $X2=1.742 $Y2=2.89
r274 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.74 $Y=2.035
+ $X2=1.74 $Y2=2.035
r275 71 79 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=0.88 $Y=2.035
+ $X2=1.74 $Y2=2.035
r276 70 75 38.6407 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=0.882 $Y=2.035
+ $X2=0.882 $Y2=2.89
r277 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.88 $Y=2.035
+ $X2=0.88 $Y2=2.035
r278 67 127 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=5.61 $Y=2.035
+ $X2=6.04 $Y2=2.035
r279 67 117 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=5.61 $Y=2.035
+ $X2=5.18 $Y2=2.035
r280 65 116 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=5.18 $Y=2.015
+ $X2=5.18 $Y2=2.035
r281 65 66 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.18 $Y=2.015
+ $X2=5.18 $Y2=1.885
r282 63 66 59.8818 $w=2.53e-07 $l=1.325e-06 $layer=LI1_cond $X=5.182 $Y=0.56
+ $X2=5.182 $Y2=1.885
r283 20 176 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=10.2
+ $Y=1.835 $X2=10.34 $Y2=2.89
r284 20 171 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=10.2
+ $Y=1.835 $X2=10.34 $Y2=2.04
r285 19 168 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=9.34
+ $Y=1.835 $X2=9.48 $Y2=2.89
r286 19 163 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=9.34
+ $Y=1.835 $X2=9.48 $Y2=2.04
r287 18 160 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=8.48
+ $Y=1.835 $X2=8.62 $Y2=2.89
r288 18 156 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=8.48
+ $Y=1.835 $X2=8.62 $Y2=2.04
r289 17 150 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=7.62
+ $Y=1.835 $X2=7.76 $Y2=2.89
r290 17 146 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.62
+ $Y=1.835 $X2=7.76 $Y2=2.04
r291 16 140 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=1.835 $X2=6.9 $Y2=2.89
r292 16 136 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=1.835 $X2=6.9 $Y2=2.04
r293 15 130 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=5.9
+ $Y=1.835 $X2=6.04 $Y2=2.89
r294 15 126 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.9
+ $Y=1.835 $X2=6.04 $Y2=2.04
r295 14 120 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.835 $X2=5.18 $Y2=2.89
r296 14 116 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.835 $X2=5.18 $Y2=2.04
r297 13 113 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=2.89
r298 13 109 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=2.04
r299 12 103 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.835 $X2=3.46 $Y2=2.89
r300 12 99 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=1.835 $X2=3.46 $Y2=2.04
r301 11 93 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.835 $X2=2.6 $Y2=2.89
r302 11 89 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.835 $X2=2.6 $Y2=2.04
r303 10 83 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.835 $X2=1.74 $Y2=2.89
r304 10 78 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.835 $X2=1.74 $Y2=2.04
r305 9 75 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.74
+ $Y=1.835 $X2=0.88 $Y2=2.89
r306 9 70 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.74
+ $Y=1.835 $X2=0.88 $Y2=2.04
r307 8 153 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.48
+ $Y=0.35 $X2=8.62 $Y2=0.56
r308 7 143 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.62
+ $Y=0.35 $X2=7.76 $Y2=0.56
r309 6 133 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.76
+ $Y=0.35 $X2=6.9 $Y2=0.56
r310 5 123 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.9
+ $Y=0.35 $X2=6.04 $Y2=0.56
r311 4 63 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.35 $X2=5.18 $Y2=0.56
r312 3 106 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.35 $X2=4.32 $Y2=0.56
r313 2 96 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.35 $X2=3.46 $Y2=0.56
r314 1 86 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.35 $X2=2.6 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_16%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 44 48
+ 52 56 60 64 67 68 70 71 72 73 75 76 78 79 81 82 83 85 103 122 123 126 129 132
r120 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r121 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r122 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r123 120 123 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r124 119 122 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r125 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r126 117 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r127 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r128 114 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.88 $Y2=0
r129 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r130 111 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.92 $Y2=0
r131 111 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r132 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r133 108 132 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=6.605 $Y=0
+ $X2=6.472 $Y2=0
r134 108 110 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.605 $Y=0
+ $X2=6.96 $Y2=0
r135 107 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r136 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r137 104 129 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.745 $Y=0
+ $X2=5.612 $Y2=0
r138 104 106 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.745 $Y=0 $X2=6
+ $Y2=0
r139 103 132 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=6.34 $Y=0
+ $X2=6.472 $Y2=0
r140 103 106 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=6
+ $Y2=0
r141 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r142 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r143 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r144 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r145 96 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r146 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r147 93 126 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.17 $Y2=0
r148 93 95 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.64 $Y2=0
r149 92 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r150 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r151 88 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=1.68 $Y2=0
r152 87 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r153 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r154 85 126 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=2.17 $Y2=0
r155 85 91 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=1.68 $Y2=0
r156 83 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r157 83 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=4.56 $Y2=0
r158 83 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r159 81 116 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=8.92 $Y=0 $X2=8.88
+ $Y2=0
r160 81 82 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.92 $Y=0 $X2=9.052
+ $Y2=0
r161 80 119 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.185 $Y=0
+ $X2=9.36 $Y2=0
r162 80 82 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=9.185 $Y=0
+ $X2=9.052 $Y2=0
r163 78 113 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.06 $Y=0 $X2=7.92
+ $Y2=0
r164 78 79 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.06 $Y=0 $X2=8.192
+ $Y2=0
r165 77 116 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.88 $Y2=0
r166 77 79 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.192 $Y2=0
r167 75 110 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.2 $Y=0 $X2=6.96
+ $Y2=0
r168 75 76 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.2 $Y=0 $X2=7.332
+ $Y2=0
r169 74 113 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=7.465 $Y=0
+ $X2=7.92 $Y2=0
r170 74 76 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=7.465 $Y=0
+ $X2=7.332 $Y2=0
r171 72 101 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.62 $Y=0 $X2=4.56
+ $Y2=0
r172 72 73 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.62 $Y=0 $X2=4.752
+ $Y2=0
r173 70 98 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.6
+ $Y2=0
r174 70 71 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.892
+ $Y2=0
r175 69 101 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=4.56 $Y2=0
r176 69 71 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=3.892 $Y2=0
r177 67 95 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.64
+ $Y2=0
r178 67 68 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.032
+ $Y2=0
r179 66 98 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.6
+ $Y2=0
r180 66 68 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.165 $Y=0
+ $X2=3.032 $Y2=0
r181 62 82 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=9.052 $Y=0.085
+ $X2=9.052 $Y2=0
r182 62 64 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=9.052 $Y=0.085
+ $X2=9.052 $Y2=0.56
r183 58 79 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=8.192 $Y=0.085
+ $X2=8.192 $Y2=0
r184 58 60 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=8.192 $Y=0.085
+ $X2=8.192 $Y2=0.56
r185 54 76 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.332 $Y=0.085
+ $X2=7.332 $Y2=0
r186 54 56 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=7.332 $Y=0.085
+ $X2=7.332 $Y2=0.56
r187 50 132 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=6.472 $Y=0.085
+ $X2=6.472 $Y2=0
r188 50 52 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=6.472 $Y=0.085
+ $X2=6.472 $Y2=0.56
r189 46 129 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.612 $Y=0.085
+ $X2=5.612 $Y2=0
r190 46 48 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=5.612 $Y=0.085
+ $X2=5.612 $Y2=0.56
r191 45 73 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.885 $Y=0
+ $X2=4.752 $Y2=0
r192 44 129 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=5.48 $Y=0
+ $X2=5.612 $Y2=0
r193 44 45 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.48 $Y=0
+ $X2=4.885 $Y2=0
r194 40 73 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.752 $Y=0.085
+ $X2=4.752 $Y2=0
r195 40 42 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=4.752 $Y=0.085
+ $X2=4.752 $Y2=0.56
r196 36 71 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.892 $Y2=0
r197 36 38 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.892 $Y2=0.56
r198 32 68 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.032 $Y=0.085
+ $X2=3.032 $Y2=0
r199 32 34 20.657 $w=2.63e-07 $l=4.75e-07 $layer=LI1_cond $X=3.032 $Y=0.085
+ $X2=3.032 $Y2=0.56
r200 28 126 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0
r201 28 30 20.2745 $w=2.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0.56
r202 9 64 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.91
+ $Y=0.35 $X2=9.05 $Y2=0.56
r203 8 60 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.05
+ $Y=0.35 $X2=8.19 $Y2=0.56
r204 7 56 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.19
+ $Y=0.35 $X2=7.33 $Y2=0.56
r205 6 52 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.35 $X2=6.47 $Y2=0.56
r206 5 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.35 $X2=5.61 $Y2=0.56
r207 4 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.61
+ $Y=0.35 $X2=4.75 $Y2=0.56
r208 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.75
+ $Y=0.35 $X2=3.89 $Y2=0.56
r209 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.35 $X2=3.03 $Y2=0.56
r210 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.35 $X2=2.17 $Y2=0.56
.ends

