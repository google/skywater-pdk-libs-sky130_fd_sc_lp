* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_562_491# D a_229_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_278_59# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1437_127# a_1406_399# a_1509_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_229_491# D a_565_59# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_2022_533# a_2064_101# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_1278_529# a_1406_399# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_229_491# a_113_63# a_312_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_312_491# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND RESET_B a_2226_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_2370_351# a_1870_127# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_1870_127# a_857_367# a_2022_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_2022_127# a_2064_101# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_229_491# a_857_367# a_1278_529# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VPWR RESET_B a_1278_529# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VGND CLK_N a_857_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_1509_127# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_857_367# a_1080_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR a_1278_529# a_1406_399# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 a_2064_101# a_1870_127# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VPWR SCE a_113_63# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 VPWR RESET_B a_2064_101# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_1406_399# a_857_367# a_1870_127# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_361_59# SCE a_229_491# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1278_529# a_1080_47# a_1364_529# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_1364_529# a_1406_399# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_2370_351# a_1870_127# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1278_529# a_857_367# a_1437_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VPWR a_2370_351# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_1870_127# a_1080_47# a_2022_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR CLK_N a_857_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VGND a_2370_351# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_229_491# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 a_1406_399# a_1080_47# a_1870_127# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X33 VPWR a_857_367# a_1080_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 VGND SCE a_113_63# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_278_59# SCD a_361_59# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_565_59# a_113_63# a_278_59# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_229_491# a_1080_47# a_1278_529# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 VPWR SCE a_562_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 a_2226_127# a_1870_127# a_2064_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
