* File: sky130_fd_sc_lp__o311ai_lp.pex.spice
* Created: Wed Sep  2 10:24:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311AI_LP%A1 3 7 9 13 14
r27 14 15 7.39264 $w=3.26e-07 $l=5e-08 $layer=POLY_cond $X=0.495 $Y=1.522
+ $X2=0.545 $Y2=1.522
r28 12 14 31.7883 $w=3.26e-07 $l=2.15e-07 $layer=POLY_cond $X=0.28 $Y=1.522
+ $X2=0.495 $Y2=1.522
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.46 $X2=0.28 $Y2=1.46
r30 9 13 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=1.46
r31 5 15 9.06345 $w=2.5e-07 $l=2.28e-07 $layer=POLY_cond $X=0.545 $Y=1.75
+ $X2=0.545 $Y2=1.522
r32 5 7 209.943 $w=2.5e-07 $l=8.45e-07 $layer=POLY_cond $X=0.545 $Y=1.75
+ $X2=0.545 $Y2=2.595
r33 1 14 20.933 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.522
r34 1 3 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%A2 3 7 9 10 11 16 17
c37 7 0 3.02941e-19 $X=1.035 $Y=2.595
r38 16 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.77
+ $X2=1.045 $Y2=1.935
r39 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.77
+ $X2=1.045 $Y2=1.605
r40 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.045
+ $Y=1.77 $X2=1.045 $Y2=1.77
r41 10 11 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.097 $Y=2.405
+ $X2=1.097 $Y2=2.775
r42 9 10 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.097 $Y=2.035
+ $X2=1.097 $Y2=2.405
r43 9 17 7.02063 $w=4.33e-07 $l=2.65e-07 $layer=LI1_cond $X=1.097 $Y=2.035
+ $X2=1.097 $Y2=1.77
r44 7 19 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.035 $Y=2.595
+ $X2=1.035 $Y2=1.935
r45 3 18 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.955 $Y=0.95
+ $X2=0.955 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%A3 1 3 8 10 11 17
r36 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=0.465 $X2=1.73 $Y2=0.465
r37 14 17 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.595 $Y=0.465
+ $X2=1.73 $Y2=0.465
r38 11 18 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=0.485
+ $X2=1.73 $Y2=0.485
r39 10 18 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=0.485 $X2=1.73
+ $Y2=0.485
r40 8 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.595 $Y=0.95 $X2=1.595
+ $Y2=1.29
r41 5 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=0.63
+ $X2=1.595 $Y2=0.465
r42 5 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.595 $Y=0.63
+ $X2=1.595 $Y2=0.95
r43 1 9 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.545 $Y=1.415
+ $X2=1.545 $Y2=1.29
r44 1 3 293.175 $w=2.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.545 $Y=1.415
+ $X2=1.545 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%B1 3 7 9 10 14
c40 14 0 1.67476e-19 $X=2.095 $Y=1.77
c41 10 0 1.74235e-19 $X=2.16 $Y=2.035
c42 3 0 1.08124e-19 $X=2.075 $Y=2.595
r43 14 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.77
+ $X2=2.095 $Y2=1.935
r44 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.77
+ $X2=2.095 $Y2=1.605
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.095
+ $Y=1.77 $X2=2.095 $Y2=1.77
r46 10 15 1.42652 $w=5.43e-07 $l=6.5e-08 $layer=LI1_cond $X=2.16 $Y=1.877
+ $X2=2.095 $Y2=1.877
r47 9 15 9.10775 $w=5.43e-07 $l=4.15e-07 $layer=LI1_cond $X=1.68 $Y=1.877
+ $X2=2.095 $Y2=1.877
r48 7 16 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.185 $Y=0.95
+ $X2=2.185 $Y2=1.605
r49 3 17 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.075 $Y=2.595
+ $X2=2.075 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%C1 3 7 9 12 13
r37 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.53
+ $X2=2.635 $Y2=1.695
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.53
+ $X2=2.635 $Y2=1.365
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.635
+ $Y=1.53 $X2=2.635 $Y2=1.53
r40 9 13 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=1.53
r41 7 15 223.608 $w=2.5e-07 $l=9e-07 $layer=POLY_cond $X=2.625 $Y=2.595
+ $X2=2.625 $Y2=1.695
r42 3 14 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=2.545 $Y=0.95
+ $X2=2.545 $Y2=1.365
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%VPWR 1 2 7 9 15 18 19 20 30 31
r42 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 22 34 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r50 22 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 20 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 20 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 18 27 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.34 $Y2=3.33
r55 17 30 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.34 $Y2=3.33
r57 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=3.245
+ $X2=2.34 $Y2=3.33
r58 13 15 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.34 $Y=3.245
+ $X2=2.34 $Y2=2.895
r59 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.24 $X2=0.28
+ $Y2=2.95
r60 7 34 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r61 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.95
r62 2 15 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=2.095 $X2=2.34 $Y2=2.895
r63 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.95
r64 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%Y 1 2 3 12 15 16 17 18 19 20 21 22 43
c48 22 0 1.08124e-19 $X=3.12 $Y=2.775
c49 15 0 1.28706e-19 $X=1.81 $Y=2.495
c50 12 0 1.67476e-19 $X=2.725 $Y=2.415
r51 44 60 1.99346 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.5 $X2=2.98
+ $Y2=2.415
r52 43 55 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=3.12 $Y=2.035 $X2=3.12
+ $Y2=2.075
r53 22 44 6.44944 $w=5.08e-07 $l=2.75e-07 $layer=LI1_cond $X=2.98 $Y=2.775
+ $X2=2.98 $Y2=2.5
r54 21 60 0.234525 $w=5.08e-07 $l=1e-08 $layer=LI1_cond $X=2.98 $Y=2.405
+ $X2=2.98 $Y2=2.415
r55 21 57 3.86967 $w=5.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.98 $Y=2.405
+ $X2=2.98 $Y2=2.24
r56 20 57 3.35371 $w=5.08e-07 $l=1.43e-07 $layer=LI1_cond $X=2.98 $Y=2.097
+ $X2=2.98 $Y2=2.24
r57 20 55 4.16556 $w=5.08e-07 $l=2.2e-08 $layer=LI1_cond $X=2.98 $Y=2.097
+ $X2=2.98 $Y2=2.075
r58 20 43 1.15244 $w=2.28e-07 $l=2.3e-08 $layer=LI1_cond $X=3.12 $Y=2.012
+ $X2=3.12 $Y2=2.035
r59 19 20 17.3869 $w=2.28e-07 $l=3.47e-07 $layer=LI1_cond $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=2.012
r60 18 19 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.665
r61 18 35 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.18
r62 17 35 4.80115 $w=2.3e-07 $l=2.3e-07 $layer=LI1_cond $X=3.12 $Y=0.95 $X2=3.12
+ $Y2=1.18
r63 17 49 9.36061 $w=4.58e-07 $l=3.6e-07 $layer=LI1_cond $X=3.12 $Y=0.95
+ $X2=2.76 $Y2=0.95
r64 17 31 4.80115 $w=2.3e-07 $l=2.3e-07 $layer=LI1_cond $X=3.12 $Y=0.95 $X2=3.12
+ $Y2=0.72
r65 16 31 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=0.555
+ $X2=3.12 $Y2=0.72
r66 13 15 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=2.415
+ $X2=1.81 $Y2=2.415
r67 12 60 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.725 $Y=2.415
+ $X2=2.98 $Y2=2.415
r68 12 13 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.725 $Y=2.415
+ $X2=1.975 $Y2=2.415
r69 3 57 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.75
+ $Y=2.095 $X2=2.89 $Y2=2.24
r70 2 15 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=1.67
+ $Y=2.095 $X2=1.81 $Y2=2.495
r71 1 49 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.74 $X2=2.76 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%VGND 1 2 7 9 13 15 17 27 28 34
r34 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r38 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r39 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r40 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r41 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r42 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 18 31 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r44 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r45 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r46 17 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.72
+ $Y2=0
r47 15 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r48 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 15 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r51 11 13 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.895
r52 7 31 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r53 7 9 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.915
r54 2 13 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.74 $X2=1.22 $Y2=0.895
r55 1 9 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.74 $X2=0.28 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_LP%A_114_148# 1 2 9 11 12 15
r31 13 15 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.89 $Y=1.255
+ $X2=1.89 $Y2=1.015
r32 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=1.34
+ $X2=1.89 $Y2=1.255
r33 11 12 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.725 $Y=1.34
+ $X2=0.875 $Y2=1.34
r34 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.75 $Y=1.255
+ $X2=0.875 $Y2=1.34
r35 7 9 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.75 $Y=1.255
+ $X2=0.75 $Y2=0.95
r36 2 15 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.74 $X2=1.89 $Y2=1.015
r37 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.74 $X2=0.71 $Y2=0.95
.ends

