* NGSPICE file created from sky130_fd_sc_lp__sdlclkp_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdlclkp_lp CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 VPWR SCE a_200_376# VPB phighvt w=1e+06u l=250000u
+  ad=1.64165e+12p pd=1.183e+07u as=2.4e+11p ps=2.48e+06u
M1001 a_1384_416# a_860_21# a_1392_192# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1002 a_698_405# a_447_376# a_93_376# VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=5.7e+11p ps=5.14e+06u
M1003 a_860_21# a_698_405# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1004 a_860_21# a_698_405# a_1016_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1005 GCLK a_1384_416# a_1548_48# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1006 a_447_376# a_356_278# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=3.9545e+11p pd=2.94e+06u as=0p ps=0u
M1007 VPWR CLK a_356_278# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1008 VPWR a_860_21# a_804_405# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1009 a_447_376# a_356_278# a_436_101# VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=8.82e+10p ps=1.26e+06u
M1010 VPWR a_860_21# a_1384_416# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1011 a_114_101# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=6.846e+11p ps=7.46e+06u
M1012 VGND CLK a_1234_192# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 a_698_405# a_356_278# a_93_376# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.373e+11p ps=2.81e+06u
M1014 a_1016_47# a_698_405# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_436_101# a_356_278# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1392_192# CLK VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1234_192# CLK a_356_278# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 a_200_376# GATE a_93_376# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_278_101# SCE a_93_376# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1020 a_1548_48# a_1384_416# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_804_405# a_356_278# a_698_405# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1022 GCLK a_1384_416# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1023 VGND SCE a_278_101# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_860_21# a_812_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 a_1384_416# CLK VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_812_47# a_447_376# a_698_405# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_93_376# GATE a_114_101# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

