* File: sky130_fd_sc_lp__sdfrbp_lp.spice
* Created: Wed Sep  2 10:34:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__sdfrbp_lp  VNB VPB SCE D SCD RESET_B CLK VPWR Q_N Q
+ VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1040 A_116_47# N_SCE_M1040_g N_A_29_47#_M1040_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_SCE_M1017_g A_116_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_342_261#_M1008_d N_SCE_M1008_g N_noxref_37_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1059 noxref_38 N_D_M1059_g N_A_342_261#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 N_noxref_39_M1004_d N_A_29_47#_M1004_g noxref_38 VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1050 N_noxref_37_M1050_d N_SCD_M1050_g N_noxref_39_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1041 N_noxref_39_M1041_d N_RESET_B_M1041_g N_VGND_M1041_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.16525 PD=1.41 PS=1.72 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_A_911_219#_M1032_d N_A_876_93#_M1032_g N_A_824_219#_M1032_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1015 N_A_342_261#_M1015_d N_A_967_193#_M1015_g N_A_911_219#_M1032_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.2724 AS=0.0588 PD=2.36 PS=0.7 NRD=169.584 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1030 A_1303_119# N_A_1147_490#_M1030_g N_A_824_219#_M1030_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_RESET_B_M1005_g A_1303_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.2753 AS=0.0504 PD=2.38 PS=0.66 NRD=171.564 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1000 A_1661_87# N_A_911_219#_M1000_g N_A_1147_490#_M1000_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1021 N_VGND_M1021_d N_A_911_219#_M1021_g A_1661_87# VNB NSHORT L=0.15 W=0.64
+ AD=0.1952 AS=0.0768 PD=1.27568 PS=0.88 NRD=46.872 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1057 A_1880_47# N_A_967_193#_M1057_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2562 PD=1.08 PS=1.67432 NRD=9.276 NRS=12.132 M=1 R=5.6
+ SA=75001.1 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_A_876_93#_M1010_d N_A_967_193#_M1010_g A_1880_47# VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1008 PD=2.25 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6
+ SA=75001.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1051 N_A_2168_439#_M1051_d N_A_876_93#_M1051_g N_A_1147_490#_M1051_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.138023 AS=0.2336 PD=1.24981 PS=2.01 NRD=0 NRS=14.988
+ M=1 R=4.26667 SA=75000.3 SB=75002 A=0.096 P=1.58 MULT=1
MM1045 A_2340_141# N_A_967_193#_M1045_g N_A_2168_439#_M1051_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0905774 PD=0.66 PS=0.820189 NRD=18.564 NRS=34.284 M=1
+ R=2.8 SA=75000.8 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_2388_115#_M1011_g A_2340_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.266725 AS=0.0504 PD=1.735 PS=0.66 NRD=34.284 NRS=18.564 M=1 R=2.8
+ SA=75001.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1054 A_2682_141# N_RESET_B_M1054_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.266725 PD=0.66 PS=1.735 NRD=18.564 NRS=222.852 M=1 R=2.8
+ SA=75002.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1035 N_A_2388_115#_M1035_d N_A_2168_439#_M1035_g A_2682_141# VNB NSHORT L=0.15
+ W=0.42 AD=0.168 AS=0.0504 PD=1.64 PS=0.66 NRD=32.856 NRS=18.564 M=1 R=2.8
+ SA=75002.9 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1026 A_3075_47# N_CLK_M1026_g N_A_967_193#_M1026_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1027 N_VGND_M1027_d N_CLK_M1027_g A_3075_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.0882 PD=1.12 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1046 A_3233_47# N_A_2168_439#_M1046_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1031 N_Q_N_M1031_d N_A_2168_439#_M1031_g A_3233_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 A_3503_137# N_A_2168_439#_M1022_g N_A_3416_137#_M1022_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_2168_439#_M1001_g A_3503_137# VNB NSHORT L=0.15 W=0.42
+ AD=0.0952 AS=0.0441 PD=0.823333 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 A_3684_53# N_A_3416_137#_M1012_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1904 PD=1.05 PS=1.64667 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1020 N_Q_M1020_d N_A_3416_137#_M1020_g A_3684_53# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1024 A_125_491# N_SCE_M1024_g N_A_29_47#_M1024_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75005.1 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_SCE_M1016_g A_125_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.184 AS=0.0672 PD=1.215 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75004.7 A=0.096 P=1.58 MULT=1
MM1013 A_342_491# N_SCE_M1013_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.184 PD=0.88 PS=1.215 NRD=19.9955 NRS=90.7973 M=1 R=4.26667
+ SA=75001.3 SB=75004 A=0.096 P=1.58 MULT=1
MM1014 N_A_342_261#_M1014_d N_D_M1014_g A_342_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.7
+ SB=75003.6 A=0.096 P=1.58 MULT=1
MM1056 A_506_491# N_A_29_47#_M1056_g N_A_342_261#_M1014_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0768 AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1023 N_VPWR_M1023_d N_SCD_M1023_g A_506_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1936 AS=0.0768 PD=1.245 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667
+ SA=75002.5 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1047 A_735_491# N_RESET_B_M1047_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1936 PD=0.88 PS=1.245 NRD=19.9955 NRS=100.037 M=1 R=4.26667
+ SA=75003.3 SB=75002 A=0.096 P=1.58 MULT=1
MM1048 N_A_342_261#_M1048_d N_RESET_B_M1048_g A_735_491# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.121419 AS=0.0768 PD=1.1834 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667
+ SA=75003.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_911_219#_M1006_d N_A_876_93#_M1006_g N_A_342_261#_M1048_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.08295 AS=0.0796811 PD=0.815 PS=0.776604 NRD=53.9386
+ NRS=30.4759 M=1 R=2.8 SA=75004.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1028 A_1020_491# N_A_967_193#_M1028_g N_A_911_219#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.18285 AS=0.08295 PD=1.275 PS=0.815 NRD=178.403 NRS=0 M=1 R=2.8
+ SA=75004.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_1147_490#_M1003_g A_1020_491# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1764 AS=0.18285 PD=1.26 PS=1.275 NRD=0 NRS=178.403 M=1 R=2.8
+ SA=75002.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1043 A_1375_535# N_RESET_B_M1043_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1764 PD=0.63 PS=1.26 NRD=23.443 NRS=262.66 M=1 R=2.8 SA=75003.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1049 N_A_911_219#_M1049_d N_RESET_B_M1049_g A_1375_535# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75004.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_1673_375# N_A_911_219#_M1002_g N_A_1147_490#_M1002_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_911_219#_M1009_g A_1673_375# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.20748 AS=0.0882 PD=1.388 PS=1.05 NRD=45.7237 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1025 A_1870_367# N_A_967_193#_M1025_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.31122 PD=1.47 PS=2.082 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_A_876_93#_M1029_d N_A_967_193#_M1029_g A_1870_367# VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1044 N_A_2168_439#_M1044_d N_A_876_93#_M1044_g N_A_2081_439#_M1044_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0952 AS=0.1197 PD=0.823333 PS=1.41 NRD=56.2829
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1042 N_A_1147_490#_M1042_d N_A_967_193#_M1042_g N_A_2168_439#_M1044_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2394 AS=0.1904 PD=2.25 PS=1.64667 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_A_2388_115#_M1018_g N_A_2081_439#_M1018_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1533 AS=0.1197 PD=1.57 PS=1.41 NRD=37.5088 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1037 N_A_2388_115#_M1037_d N_A_2168_439#_M1037_g N_A_2523_397#_M1037_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.138912 AS=0.1197 PD=1.42 PS=1.41 NRD=129.331 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 A_2719_518# N_RESET_B_M1038_g N_A_2388_115#_M1037_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.138912 PD=0.63 PS=1.42 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_RESET_B_M1036_g A_2719_518# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_A_2523_397#_M1019_d N_A_2168_439#_M1019_g N_VPWR_M1036_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1052 A_3075_357# N_CLK_M1052_g N_A_967_193#_M1052_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3591 PD=1.47 PS=3.09 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1055 N_VPWR_M1055_d N_CLK_M1055_g A_3075_357# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75001 A=0.189 P=2.82 MULT=1
MM1033 A_3233_357# N_A_2168_439#_M1033_g N_VPWR_M1055_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1007 N_Q_N_M1007_d N_A_2168_439#_M1007_g A_3233_357# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1034 A_3503_367# N_A_2168_439#_M1034_g N_A_3416_137#_M1034_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=15.3857 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1039 N_VPWR_M1039_d N_A_2168_439#_M1039_g A_3503_367# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.144674 AS=0.0672 PD=1.11495 PS=0.85 NRD=36.1495 NRS=15.3857 M=1
+ R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1053 A_3684_367# N_A_3416_137#_M1053_g N_VPWR_M1039_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1323 AS=0.284826 PD=1.47 PS=2.19505 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1058 N_Q_M1058_d N_A_3416_137#_M1058_g A_3684_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX60_noxref VNB VPB NWDIODE A=33.6584 P=44.23
c_378 VPB 0 1.20402e-19 $X=0 $Y=3.085
c_2972 A_1303_119# 0 1.97601e-20 $X=6.515 $Y=0.595
*
.include "sky130_fd_sc_lp__sdfrbp_lp.pxi.spice"
*
.ends
*
*
