* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and3b_2 A_N B C VGND VNB VPB VPWR X
M1000 a_204_27# C VPWR VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.0983e+12p ps=8.79e+06u
M1001 VPWR a_204_27# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1002 a_204_27# a_27_137# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_489_137# C VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.729e+11p ps=6.17e+06u
M1004 VPWR B a_204_27# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A_N a_27_137# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 a_561_137# B a_489_137# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1007 a_204_27# a_27_137# a_561_137# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1008 VPWR A_N a_27_137# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 X a_204_27# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1010 VGND a_204_27# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_204_27# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
