* File: sky130_fd_sc_lp__o41a_lp.spice
* Created: Wed Sep  2 10:27:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o41a_lp  VNB VPB A1 A2 A3 A4 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A1_M1002_g N_A_31_57#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1197 PD=0.86 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_31_57#_M1003_d N_A2_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.0924 PD=0.735 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A3_M1000_g N_A_31_57#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.06615 PD=0.745 PS=0.735 NRD=12.852 NRS=9.996 M=1 R=2.8
+ SA=75001.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_A_31_57#_M1009_d N_A4_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.06825 PD=0.7 PS=0.745 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_457_412#_M1011_d N_B1_M1011_g N_A_31_57#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_708_47# N_A_457_412#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_457_412#_M1001_g A_708_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_137_412# N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1010 A_235_412# N_A2_M1010_g A_137_412# VPB PHIGHVT L=0.25 W=1 AD=0.16 AS=0.12
+ PD=1.32 PS=1.24 NRD=20.6653 NRS=12.7853 M=1 R=4 SA=125001 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1007 A_349_412# N_A3_M1007_g A_235_412# VPB PHIGHVT L=0.25 W=1 AD=0.145
+ AS=0.16 PD=1.29 PS=1.32 NRD=17.7103 NRS=20.6653 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1004 N_A_457_412#_M1004_d N_A4_M1004_g A_349_412# VPB PHIGHVT L=0.25 W=1
+ AD=0.2825 AS=0.145 PD=1.565 PS=1.29 NRD=56.145 NRS=17.7103 M=1 R=4 SA=125002
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_B1_M1012_g N_A_457_412#_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1975 AS=0.2825 PD=1.395 PS=1.565 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1005 N_X_M1005_d N_A_457_412#_M1005_g N_VPWR_M1012_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1975 PD=2.57 PS=1.395 NRD=0 NRS=22.6353 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o41a_lp.pxi.spice"
*
.ends
*
*
