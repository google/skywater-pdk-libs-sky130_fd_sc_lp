* File: sky130_fd_sc_lp__nor2_2.pex.spice
* Created: Wed Sep  2 10:07:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_2%A 1 3 6 8 10 13 15 16 24
r43 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.48 $Y=1.375
+ $X2=0.91 $Y2=1.375
r44 20 23 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.345 $Y=1.375
+ $X2=0.48 $Y2=1.375
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.345
+ $Y=1.375 $X2=0.345 $Y2=1.375
r46 16 21 9.6872 $w=3.43e-07 $l=2.9e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=1.375
r47 15 21 2.67233 $w=3.43e-07 $l=8e-08 $layer=LI1_cond $X=0.257 $Y=1.295
+ $X2=0.257 $Y2=1.375
r48 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.54
+ $X2=0.91 $Y2=1.375
r49 11 13 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.91 $Y=1.54
+ $X2=0.91 $Y2=2.465
r50 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.21
+ $X2=0.91 $Y2=1.375
r51 8 10 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.91 $Y=1.21
+ $X2=0.91 $Y2=0.665
r52 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.54
+ $X2=0.48 $Y2=1.375
r53 4 6 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.48 $Y=1.54 $X2=0.48
+ $Y2=2.465
r54 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.21
+ $X2=0.48 $Y2=1.375
r55 1 3 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.48 $Y=1.21 $X2=0.48
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_2%B 3 7 11 15 17 18 25 26
c50 26 0 9.26868e-20 $X=1.77 $Y=1.51
r51 24 26 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.36 $Y=1.51
+ $X2=1.77 $Y2=1.51
r52 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.36
+ $Y=1.51 $X2=1.36 $Y2=1.51
r53 21 24 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.34 $Y=1.51 $X2=1.36
+ $Y2=1.51
r54 18 25 5.67357 $w=3.23e-07 $l=1.6e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.36 $Y2=1.587
r55 17 18 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=1.2 $Y2=1.587
r56 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.675
+ $X2=1.77 $Y2=1.51
r57 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.77 $Y=1.675
+ $X2=1.77 $Y2=2.465
r58 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.345
+ $X2=1.77 $Y2=1.51
r59 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.77 $Y=1.345
+ $X2=1.77 $Y2=0.665
r60 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.675
+ $X2=1.34 $Y2=1.51
r61 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.34 $Y=1.675 $X2=1.34
+ $Y2=2.465
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.345
+ $X2=1.34 $Y2=1.51
r63 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.34 $Y=1.345 $X2=1.34
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_2%A_28_367# 1 2 3 10 12 14 16 17 18 20 22
c32 16 0 9.26868e-20 $X=1.12 $Y=2.09
r33 20 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.905
+ $X2=2.17 $Y2=2.99
r34 20 22 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=2.17 $Y=2.905
+ $X2=2.17 $Y2=1.985
r35 19 29 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.21 $Y=2.99 $X2=1.12
+ $Y2=2.99
r36 18 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=2.17 $Y2=2.99
r37 18 19 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=1.21 $Y2=2.99
r38 17 29 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.905
+ $X2=1.12 $Y2=2.99
r39 16 27 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.09 $X2=1.12
+ $Y2=2.005
r40 16 17 50.2172 $w=1.78e-07 $l=8.15e-07 $layer=LI1_cond $X=1.12 $Y=2.09
+ $X2=1.12 $Y2=2.905
r41 15 25 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.36 $Y=2.005
+ $X2=0.23 $Y2=2.005
r42 14 27 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.03 $Y=2.005 $X2=1.12
+ $Y2=2.005
r43 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.03 $Y=2.005
+ $X2=0.36 $Y2=2.005
r44 10 25 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.09 $X2=0.23
+ $Y2=2.005
r45 10 12 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.23 $Y=2.09
+ $X2=0.23 $Y2=2.91
r46 3 31 400 $w=1.7e-07 $l=1.20913e-06 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.835 $X2=2.13 $Y2=2.91
r47 3 22 400 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.835 $X2=2.13 $Y2=1.985
r48 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.91
r49 2 27 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.085
r50 1 25 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.085
r51 1 12 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_2%VPWR 1 6 8 10 20 21 24
r31 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r34 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=3.33
+ $X2=0.695 $Y2=3.33
r35 15 17 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.695 $Y2=3.33
r39 10 12 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 8 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r41 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.72
+ $Y2=3.33
r42 8 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r44 4 6 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.385
r45 1 6 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_2%Y 1 2 3 12 14 15 21 22 25 26 27 31
r41 26 27 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.612 $Y=0.555
+ $X2=1.612 $Y2=0.925
r42 26 31 5.10098 $w=3.03e-07 $l=1.35e-07 $layer=LI1_cond $X=1.612 $Y=0.555
+ $X2=1.612 $Y2=0.42
r43 24 27 5.66775 $w=3.03e-07 $l=1.5e-07 $layer=LI1_cond $X=1.612 $Y=1.075
+ $X2=1.612 $Y2=0.925
r44 24 25 3.80849 $w=2.42e-07 $l=1.14237e-07 $layer=LI1_cond $X=1.612 $Y=1.075
+ $X2=1.667 $Y2=1.165
r45 21 22 8.12202 $w=4.93e-07 $l=1.25e-07 $layer=LI1_cond $X=1.627 $Y=2.045
+ $X2=1.627 $Y2=1.92
r46 18 25 3.80849 $w=2.42e-07 $l=1.56665e-07 $layer=LI1_cond $X=1.785 $Y=1.255
+ $X2=1.667 $Y2=1.165
r47 18 22 40.9747 $w=1.78e-07 $l=6.65e-07 $layer=LI1_cond $X=1.785 $Y=1.255
+ $X2=1.785 $Y2=1.92
r48 14 25 2.64776 $w=1.7e-07 $l=2.09485e-07 $layer=LI1_cond $X=1.46 $Y=1.17
+ $X2=1.667 $Y2=1.165
r49 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.46 $Y=1.17
+ $X2=0.79 $Y2=1.17
r50 10 15 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.7 $Y=1.085
+ $X2=0.79 $Y2=1.17
r51 10 12 40.9747 $w=1.78e-07 $l=6.65e-07 $layer=LI1_cond $X=0.7 $Y=1.085
+ $X2=0.7 $Y2=0.42
r52 3 21 300 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.835 $X2=1.555 $Y2=2.045
r53 2 31 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.415
+ $Y=0.245 $X2=1.555 $Y2=0.42
r54 1 12 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.245 $X2=0.695 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_2%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
r34 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 33 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r37 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r38 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.125
+ $Y2=0
r39 30 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.68
+ $Y2=0
r40 29 41 3.90852 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.167
+ $Y2=0
r41 29 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.68
+ $Y2=0
r42 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r43 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 25 35 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r45 25 27 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r46 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.125
+ $Y2=0
r47 24 27 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r48 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r49 22 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r50 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 18 41 3.23464 $w=2.5e-07 $l=1.43332e-07 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.167 $Y2=0
r52 18 20 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=2.06 $Y=0.085
+ $X2=2.06 $Y2=0.39
r53 14 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0
r54 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0.39
r55 10 35 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.215 $Y2=0
r56 10 12 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.39
r57 3 20 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=1.845
+ $Y=0.245 $X2=2.02 $Y2=0.39
r58 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.245 $X2=1.125 $Y2=0.39
r59 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.245 $X2=0.265 $Y2=0.39
.ends

