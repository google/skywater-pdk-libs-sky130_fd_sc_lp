* File: sky130_fd_sc_lp__einvp_1.pxi.spice
* Created: Fri Aug 28 10:33:44 2020
* 
x_PM_SKY130_FD_SC_LP__EINVP_1%A N_A_M1003_g N_A_M1005_g A A N_A_c_43_n
+ PM_SKY130_FD_SC_LP__EINVP_1%A
x_PM_SKY130_FD_SC_LP__EINVP_1%A_207_302# N_A_207_302#_M1004_d
+ N_A_207_302#_M1000_d N_A_207_302#_M1002_g N_A_207_302#_c_73_n
+ N_A_207_302#_c_74_n N_A_207_302#_c_75_n N_A_207_302#_c_69_n
+ N_A_207_302#_c_70_n N_A_207_302#_c_71_n PM_SKY130_FD_SC_LP__EINVP_1%A_207_302#
x_PM_SKY130_FD_SC_LP__EINVP_1%TE N_TE_c_110_n N_TE_M1001_g N_TE_c_111_n
+ N_TE_M1000_g N_TE_c_113_n N_TE_M1004_g TE TE N_TE_c_114_n N_TE_c_115_n
+ N_TE_c_116_n PM_SKY130_FD_SC_LP__EINVP_1%TE
x_PM_SKY130_FD_SC_LP__EINVP_1%Z N_Z_M1003_s N_Z_M1005_s Z Z Z Z Z Z Z
+ N_Z_c_153_n Z PM_SKY130_FD_SC_LP__EINVP_1%Z
x_PM_SKY130_FD_SC_LP__EINVP_1%VPWR N_VPWR_M1002_d N_VPWR_c_185_n VPWR
+ N_VPWR_c_186_n N_VPWR_c_187_n N_VPWR_c_184_n N_VPWR_c_189_n
+ PM_SKY130_FD_SC_LP__EINVP_1%VPWR
x_PM_SKY130_FD_SC_LP__EINVP_1%VGND N_VGND_M1001_d N_VGND_c_207_n VGND
+ N_VGND_c_208_n N_VGND_c_209_n N_VGND_c_210_n N_VGND_c_211_n
+ PM_SKY130_FD_SC_LP__EINVP_1%VGND
cc_1 VNB N_A_M1003_g 0.0273032f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.655
cc_2 VNB A 0.0238152f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_43_n 0.0491511f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.51
cc_4 VNB N_A_207_302#_c_69_n 0.0460564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_207_302#_c_70_n 0.0147085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_207_302#_c_71_n 0.0016919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_TE_c_110_n 0.0190917f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.295
cc_8 VNB N_TE_c_111_n 0.0133965f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.725
cc_9 VNB N_TE_M1000_g 0.00778268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_TE_c_113_n 0.0645293f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_TE_c_114_n 0.0280166f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_12 VNB N_TE_c_115_n 0.00480239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_TE_c_116_n 9.1847e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB Z 0.00847297f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_Z_c_153_n 0.0336819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_184_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_207_n 0.0255979f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.5
cc_18 VNB N_VGND_c_208_n 0.02848f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.46
cc_19 VNB N_VGND_c_209_n 0.0193537f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_20 VNB N_VGND_c_210_n 0.160525f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_21 VNB N_VGND_c_211_n 0.0151955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A_M1005_g 0.0288185f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.5
cc_23 VPB A 0.0170522f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_24 VPB N_A_c_43_n 0.0197875f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.51
cc_25 VPB N_A_207_302#_M1002_g 0.021284f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_26 VPB N_A_207_302#_c_73_n 0.00392358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_A_207_302#_c_74_n 0.0349135f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.46
cc_28 VPB N_A_207_302#_c_75_n 0.0231939f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.725
cc_29 VPB N_A_207_302#_c_69_n 0.00245284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_A_207_302#_c_70_n 0.0155678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_207_302#_c_71_n 0.00369155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_TE_M1000_g 0.0372418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB Z 0.00718079f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB Z 0.0361861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB Z 0.0135833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_185_n 0.0281033f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.5
cc_37 VPB N_VPWR_c_186_n 0.0341284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_187_n 0.0298284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_184_n 0.0925774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_189_n 0.00659812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 N_A_M1005_g N_A_207_302#_M1002_g 0.0418292f $X=0.73 $Y=2.5 $X2=0 $Y2=0
cc_42 N_A_c_43_n N_A_207_302#_c_70_n 0.0435802f $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_43 N_A_c_43_n N_A_207_302#_c_71_n 3.34714e-19 $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_44 N_A_M1003_g N_TE_c_110_n 0.0304052f $X=0.565 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_45 N_A_c_43_n N_TE_c_111_n 0.0304052f $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_46 N_A_c_43_n N_TE_c_115_n 4.1248e-19 $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_47 N_A_M1003_g Z 0.00788445f $X=0.565 $Y=0.655 $X2=0 $Y2=0
cc_48 N_A_M1005_g Z 0.00798549f $X=0.73 $Y=2.5 $X2=0 $Y2=0
cc_49 A Z 0.0437169f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A_c_43_n Z 0.0190042f $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_51 N_A_M1005_g Z 0.0165028f $X=0.73 $Y=2.5 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_Z_c_153_n 0.0288258f $X=0.565 $Y=0.655 $X2=0 $Y2=0
cc_53 A N_Z_c_153_n 0.0234623f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A_c_43_n N_Z_c_153_n 0.00152468f $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_55 N_A_M1005_g Z 0.00533228f $X=0.73 $Y=2.5 $X2=0 $Y2=0
cc_56 A Z 0.00953554f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A_c_43_n Z 0.00831013f $X=0.565 $Y=1.51 $X2=0 $Y2=0
cc_58 N_A_M1005_g N_VPWR_c_185_n 0.00157658f $X=0.73 $Y=2.5 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_VPWR_c_186_n 0.00305149f $X=0.73 $Y=2.5 $X2=0 $Y2=0
cc_60 N_A_M1005_g N_VPWR_c_184_n 0.00461254f $X=0.73 $Y=2.5 $X2=0 $Y2=0
cc_61 N_A_M1003_g N_VGND_c_208_n 0.00357668f $X=0.565 $Y=0.655 $X2=0 $Y2=0
cc_62 N_A_M1003_g N_VGND_c_210_n 0.00627715f $X=0.565 $Y=0.655 $X2=0 $Y2=0
cc_63 N_A_207_302#_M1002_g N_TE_M1000_g 0.0112395f $X=1.11 $Y=2.5 $X2=0 $Y2=0
cc_64 N_A_207_302#_c_73_n N_TE_M1000_g 0.0110706f $X=1.7 $Y=1.775 $X2=0 $Y2=0
cc_65 N_A_207_302#_c_74_n N_TE_M1000_g 0.0118851f $X=1.865 $Y=2.215 $X2=0 $Y2=0
cc_66 N_A_207_302#_c_75_n N_TE_M1000_g 0.00491772f $X=2.135 $Y=1.685 $X2=0 $Y2=0
cc_67 N_A_207_302#_c_69_n N_TE_M1000_g 0.00410716f $X=2.11 $Y=0.865 $X2=0 $Y2=0
cc_68 N_A_207_302#_c_71_n N_TE_M1000_g 0.00129564f $X=1.415 $Y=1.712 $X2=0 $Y2=0
cc_69 N_A_207_302#_c_75_n N_TE_c_113_n 0.00595023f $X=2.135 $Y=1.685 $X2=0 $Y2=0
cc_70 N_A_207_302#_c_69_n N_TE_c_113_n 0.0143957f $X=2.11 $Y=0.865 $X2=0 $Y2=0
cc_71 N_A_207_302#_c_70_n N_TE_c_113_n 0.0207635f $X=1.2 $Y=1.675 $X2=0 $Y2=0
cc_72 N_A_207_302#_c_73_n N_TE_c_114_n 8.48566e-19 $X=1.7 $Y=1.775 $X2=0 $Y2=0
cc_73 N_A_207_302#_c_70_n N_TE_c_114_n 0.0210769f $X=1.2 $Y=1.675 $X2=0 $Y2=0
cc_74 N_A_207_302#_c_71_n N_TE_c_114_n 6.52345e-19 $X=1.415 $Y=1.712 $X2=0 $Y2=0
cc_75 N_A_207_302#_c_73_n N_TE_c_115_n 0.00880845f $X=1.7 $Y=1.775 $X2=0 $Y2=0
cc_76 N_A_207_302#_c_70_n N_TE_c_115_n 0.00199748f $X=1.2 $Y=1.675 $X2=0 $Y2=0
cc_77 N_A_207_302#_c_71_n N_TE_c_115_n 0.0282981f $X=1.415 $Y=1.712 $X2=0 $Y2=0
cc_78 N_A_207_302#_c_73_n N_TE_c_116_n 0.0175162f $X=1.7 $Y=1.775 $X2=0 $Y2=0
cc_79 N_A_207_302#_c_69_n N_TE_c_116_n 0.0255666f $X=2.11 $Y=0.865 $X2=0 $Y2=0
cc_80 N_A_207_302#_M1002_g Z 0.0116916f $X=1.11 $Y=2.5 $X2=0 $Y2=0
cc_81 N_A_207_302#_c_70_n Z 0.00219925f $X=1.2 $Y=1.675 $X2=0 $Y2=0
cc_82 N_A_207_302#_c_71_n Z 0.0243454f $X=1.415 $Y=1.712 $X2=0 $Y2=0
cc_83 N_A_207_302#_M1002_g N_VPWR_c_185_n 0.0181221f $X=1.11 $Y=2.5 $X2=0 $Y2=0
cc_84 N_A_207_302#_c_74_n N_VPWR_c_185_n 0.0148031f $X=1.865 $Y=2.215 $X2=0
+ $Y2=0
cc_85 N_A_207_302#_c_70_n N_VPWR_c_185_n 0.00116678f $X=1.2 $Y=1.675 $X2=0 $Y2=0
cc_86 N_A_207_302#_c_71_n N_VPWR_c_185_n 0.0280617f $X=1.415 $Y=1.712 $X2=0
+ $Y2=0
cc_87 N_A_207_302#_M1002_g N_VPWR_c_186_n 0.00411131f $X=1.11 $Y=2.5 $X2=0 $Y2=0
cc_88 N_A_207_302#_M1002_g N_VPWR_c_184_n 0.00780741f $X=1.11 $Y=2.5 $X2=0 $Y2=0
cc_89 N_A_207_302#_c_69_n N_VGND_c_209_n 0.00462376f $X=2.11 $Y=0.865 $X2=0
+ $Y2=0
cc_90 N_A_207_302#_c_69_n N_VGND_c_210_n 0.00804028f $X=2.11 $Y=0.865 $X2=0
+ $Y2=0
cc_91 N_TE_c_110_n Z 0.00725997f $X=0.955 $Y=1.15 $X2=0 $Y2=0
cc_92 N_TE_c_115_n Z 0.0164268f $X=1.585 $Y=1.285 $X2=0 $Y2=0
cc_93 N_TE_M1000_g N_VPWR_c_185_n 0.00592578f $X=1.65 $Y=2.21 $X2=0 $Y2=0
cc_94 N_TE_M1000_g N_VPWR_c_187_n 0.00292498f $X=1.65 $Y=2.21 $X2=0 $Y2=0
cc_95 N_TE_M1000_g N_VPWR_c_184_n 0.00397372f $X=1.65 $Y=2.21 $X2=0 $Y2=0
cc_96 N_TE_c_110_n N_VGND_c_207_n 0.0067928f $X=0.955 $Y=1.15 $X2=0 $Y2=0
cc_97 N_TE_c_113_n N_VGND_c_207_n 0.0160464f $X=1.875 $Y=1.15 $X2=0 $Y2=0
cc_98 N_TE_c_114_n N_VGND_c_207_n 0.0132218f $X=1.575 $Y=1.332 $X2=0 $Y2=0
cc_99 N_TE_c_115_n N_VGND_c_207_n 0.04131f $X=1.585 $Y=1.285 $X2=0 $Y2=0
cc_100 N_TE_c_116_n N_VGND_c_207_n 0.0170955f $X=1.705 $Y=1.285 $X2=0 $Y2=0
cc_101 N_TE_c_110_n N_VGND_c_208_n 0.00585385f $X=0.955 $Y=1.15 $X2=0 $Y2=0
cc_102 N_TE_c_113_n N_VGND_c_209_n 0.00332367f $X=1.875 $Y=1.15 $X2=0 $Y2=0
cc_103 N_TE_c_110_n N_VGND_c_210_n 0.011835f $X=0.955 $Y=1.15 $X2=0 $Y2=0
cc_104 N_TE_c_113_n N_VGND_c_210_n 0.00387424f $X=1.875 $Y=1.15 $X2=0 $Y2=0
cc_105 Z A_161_400# 0.00848007f $X=0.635 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_106 Z A_161_400# 0.00243763f $X=0.72 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_107 Z N_VPWR_c_185_n 0.0534473f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_108 Z N_VPWR_c_186_n 0.0295963f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_109 Z N_VPWR_c_184_n 0.0188987f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_110 N_Z_c_153_n A_128_47# 0.00136237f $X=0.35 $Y=0.38 $X2=-0.19 $Y2=-0.245
cc_111 N_Z_c_153_n N_VGND_c_208_n 0.0419729f $X=0.35 $Y=0.38 $X2=0 $Y2=0
cc_112 N_Z_M1003_s N_VGND_c_210_n 0.00215158f $X=0.225 $Y=0.235 $X2=0 $Y2=0
cc_113 N_Z_c_153_n N_VGND_c_210_n 0.0255996f $X=0.35 $Y=0.38 $X2=0 $Y2=0
cc_114 A_128_47# N_VGND_c_210_n 0.00248661f $X=0.64 $Y=0.235 $X2=0.745 $Y2=1.04
