* File: sky130_fd_sc_lp__nor2_1.spice
* Created: Wed Sep  2 10:07:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor2_1.pex.spice"
.subckt sky130_fd_sc_lp__nor2_1  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1000 A_116_367# N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26 AD=0.1512
+ AS=0.3339 PD=1.5 PS=3.05 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g A_116_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.3339
+ AS=0.1512 PD=3.05 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
c_94 A_116_367# 0 6.79148e-20 $X=0.58 $Y=1.835
*
.include "sky130_fd_sc_lp__nor2_1.pxi.spice"
*
.ends
*
*
