* File: sky130_fd_sc_lp__maj3_2.spice
* Created: Fri Aug 28 10:43:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__maj3_2.pex.spice"
.subckt sky130_fd_sc_lp__maj3_2  VNB VPB C A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C	C
* VPB	VPB
* VNB	VNB
MM1002 A_154_49# N_C_M1002_g N_A_59_491#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g A_154_49# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75002.9
+ A=0.063 P=1.14 MULT=1
MM1006 A_318_49# N_A_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_59_491#_M1007_d N_B_M1007_g A_318_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1014 A_482_49# N_B_M1014_g N_A_59_491#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_C_M1015_g A_482_49# VNB NSHORT L=0.15 W=0.42 AD=0.0854
+ AS=0.0504 PD=0.8 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_59_491#_M1001_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1708 PD=1.12 PS=1.6 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.5
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1012 N_X_M1001_d N_A_59_491#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3738 PD=1.12 PS=2.57 NRD=0 NRS=22.848 M=1 R=5.6 SA=75001.9
+ SB=75000.4 A=0.126 P=1.98 MULT=1
MM1008 A_146_491# N_C_M1008_g N_A_59_491#_M1008_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g A_146_491# VPB PHIGHVT L=0.15 W=0.64 AD=0.0896
+ AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.6 SB=75003
+ A=0.096 P=1.58 MULT=1
MM1000 A_310_491# N_A_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75001 SB=75002.6
+ A=0.096 P=1.58 MULT=1
MM1010 N_A_59_491#_M1010_d N_B_M1010_g A_310_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.4
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 A_474_491# N_B_M1004_g N_A_59_491#_M1010_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_C_M1011_g A_474_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.172935 AS=0.0768 PD=1.22611 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667
+ SA=75002.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1011_d N_A_59_491#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.340465 AS=0.1764 PD=2.41389 PS=1.54 NRD=43.7734 NRS=0 M=1 R=8.4
+ SA=75001.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_59_491#_M1013_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__maj3_2.pxi.spice"
*
.ends
*
*
