* File: sky130_fd_sc_lp__o211ai_1.pex.spice
* Created: Fri Aug 28 11:02:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211AI_1%A1 3 7 9 10 17
c28 9 0 1.85267e-19 $X=0.24 $Y=1.295
r29 14 17 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.375
+ $X2=0.475 $Y2=1.375
r30 9 10 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295 $X2=0.26
+ $Y2=1.665
r31 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.375 $X2=0.27 $Y2=1.375
r32 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=1.375
r33 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=2.465
r34 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.21
+ $X2=0.475 $Y2=1.375
r35 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.475 $Y=1.21
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_1%A2 3 7 8 9 10 11 12 19 20 21
c46 19 0 1.73662e-19 $X=0.925 $Y=1.35
c47 3 0 1.85267e-19 $X=0.835 $Y=2.465
r48 23 36 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.515
+ $X2=0.725 $Y2=1.35
r49 20 36 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.925 $Y=1.35 $X2=0.725
+ $Y2=1.35
r50 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.515
r51 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.185
r52 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.35 $X2=0.925 $Y2=1.35
r53 11 12 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=2.405
+ $X2=0.725 $Y2=2.775
r54 10 11 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=2.035
+ $X2=0.725 $Y2=2.405
r55 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=2.035
r56 9 23 7.20277 $w=2.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=1.515
r57 8 36 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.72 $Y=1.35 $X2=0.725
+ $Y2=1.35
r58 7 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.015 $Y=0.655
+ $X2=1.015 $Y2=1.185
r59 3 22 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.835 $Y=2.465
+ $X2=0.835 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_1%B1 3 6 8 9 10 11 18 21 30
c46 21 0 3.68135e-20 $X=1.465 $Y=1.725
c47 8 0 1.73662e-19 $X=1.68 $Y=0.555
r48 30 32 2.56098 $w=2.23e-07 $l=5e-08 $layer=LI1_cond $X=1.682 $Y=1.295
+ $X2=1.682 $Y2=1.345
r49 18 21 54.9546 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.465 $Y=1.51
+ $X2=1.465 $Y2=1.725
r50 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.51
+ $X2=1.465 $Y2=1.345
r51 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.51 $X2=1.465 $Y2=1.51
r52 11 19 3.7453 $w=4.93e-07 $l=1.55e-07 $layer=LI1_cond $X=1.547 $Y=1.665
+ $X2=1.547 $Y2=1.51
r53 10 19 3.57615 $w=4.93e-07 $l=1.48e-07 $layer=LI1_cond $X=1.547 $Y=1.362
+ $X2=1.547 $Y2=1.51
r54 10 32 4.00898 $w=4.93e-07 $l=1.7e-08 $layer=LI1_cond $X=1.547 $Y=1.362
+ $X2=1.547 $Y2=1.345
r55 10 30 0.921954 $w=2.23e-07 $l=1.8e-08 $layer=LI1_cond $X=1.682 $Y=1.277
+ $X2=1.682 $Y2=1.295
r56 9 10 18.0293 $w=2.23e-07 $l=3.52e-07 $layer=LI1_cond $X=1.682 $Y=0.925
+ $X2=1.682 $Y2=1.277
r57 8 9 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.682 $Y=0.555
+ $X2=1.682 $Y2=0.925
r58 6 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.555 $Y=0.655
+ $X2=1.555 $Y2=1.345
r59 3 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.375 $Y=2.465
+ $X2=1.375 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_1%C1 3 7 9 14 15
c31 15 0 3.68135e-20 $X=2.1 $Y=1.46
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.1
+ $Y=1.46 $X2=2.1 $Y2=1.46
r33 11 14 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.915 $Y=1.46
+ $X2=2.1 $Y2=1.46
r34 9 15 7.05226 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=2.132 $Y=1.665
+ $X2=2.132 $Y2=1.46
r35 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.625
+ $X2=1.915 $Y2=1.46
r36 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.915 $Y=1.625
+ $X2=1.915 $Y2=2.465
r37 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.295
+ $X2=1.915 $Y2=1.46
r38 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.915 $Y=1.295
+ $X2=1.915 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_1%VPWR 1 2 7 9 15 17 19 26 27 33
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.645 $Y2=3.33
r39 24 26 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 23 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 20 30 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r43 20 22 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=3.33
+ $X2=1.645 $Y2=3.33
r45 19 22 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.48 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 17 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 17 23 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=3.33
r49 13 15 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=2.39
r50 9 12 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.26 $Y=2.005
+ $X2=0.26 $Y2=2.95
r51 7 30 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r52 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r53 2 15 300 $w=1.7e-07 $l=6.45174e-07 $layer=licon1_PDIFF $count=2 $X=1.45
+ $Y=1.835 $X2=1.645 $Y2=2.39
r54 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r55 1 9 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_1%Y 1 2 3 10 12 14 18 19 20 21 22 23 24 51
r44 24 46 4.56005 $w=7.98e-07 $l=3.05e-07 $layer=LI1_cond $X=2.38 $Y=2.775
+ $X2=2.38 $Y2=2.47
r45 23 46 0.971814 $w=7.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.38 $Y=2.405
+ $X2=2.38 $Y2=2.47
r46 22 23 3.99536 $w=9.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.38 $Y=2.12
+ $X2=2.38 $Y2=2.405
r47 21 22 8.5987 $w=4.78e-07 $l=2.85e-07 $layer=LI1_cond $X=2.625 $Y=1.665
+ $X2=2.625 $Y2=1.95
r48 20 21 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=1.295
+ $X2=2.625 $Y2=1.665
r49 20 57 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=2.625 $Y=1.295
+ $X2=2.625 $Y2=1.095
r50 19 57 7.2865 $w=8.13e-07 $l=1.7e-07 $layer=LI1_cond $X=2.372 $Y=0.925
+ $X2=2.372 $Y2=1.095
r51 18 19 5.43005 $w=8.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.372 $Y=0.555
+ $X2=2.372 $Y2=0.925
r52 18 51 2.56827 $w=8.13e-07 $l=1.75e-07 $layer=LI1_cond $X=2.372 $Y=0.555
+ $X2=2.372 $Y2=0.38
r53 15 17 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.28 $Y=2.035
+ $X2=1.147 $Y2=2.035
r54 14 22 5.8014 $w=1.7e-07 $l=4e-07 $layer=LI1_cond $X=1.98 $Y=2.035 $X2=2.38
+ $Y2=2.035
r55 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.98 $Y=2.035 $X2=1.28
+ $Y2=2.035
r56 10 17 2.82608 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.147 $Y=2.12
+ $X2=1.147 $Y2=2.035
r57 10 12 34.3558 $w=2.63e-07 $l=7.9e-07 $layer=LI1_cond $X=1.147 $Y=2.12
+ $X2=1.147 $Y2=2.91
r58 3 22 300 $w=1.7e-07 $l=5.71314e-07 $layer=licon1_PDIFF $count=2 $X=1.99
+ $Y=1.835 $X2=2.47 $Y2=2.035
r59 3 46 150 $w=1.7e-07 $l=8.41442e-07 $layer=licon1_PDIFF $count=4 $X=1.99
+ $Y=1.835 $X2=2.47 $Y2=2.47
r60 2 17 400 $w=1.7e-07 $l=3.68511e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=1.835 $X2=1.115 $Y2=2.115
r61 2 12 400 $w=1.7e-07 $l=1.17303e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=1.835 $X2=1.115 $Y2=2.91
r62 1 51 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=1.99
+ $Y=0.235 $X2=2.47 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_1%A_27_47# 1 2 9 11 12 15
r27 13 15 17.8105 $w=2.73e-07 $l=4.25e-07 $layer=LI1_cond $X=1.262 $Y=0.845
+ $X2=1.262 $Y2=0.42
r28 11 13 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=1.125 $Y=0.93
+ $X2=1.262 $Y2=0.845
r29 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.125 $Y=0.93
+ $X2=0.425 $Y2=0.93
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.845
+ $X2=0.425 $Y2=0.93
r31 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.26 $Y=0.845 $X2=0.26
+ $Y2=0.38
r32 2 15 91 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.235 $X2=1.29 $Y2=0.42
r33 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_1%VGND 1 6 8 10 20 21 24
r30 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r32 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r33 17 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r34 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.76
+ $Y2=0
r36 15 17 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.2
+ $Y2=0
r37 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r38 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.76
+ $Y2=0
r40 10 12 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.24
+ $Y2=0
r41 8 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r42 8 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r43 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0
r44 4 6 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.76 $Y=0.085 $X2=0.76
+ $Y2=0.55
r45 1 6 182 $w=1.7e-07 $l=4.06663e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.76 $Y2=0.55
.ends

