* File: sky130_fd_sc_lp__mux2_lp.pex.spice
* Created: Wed Sep  2 10:00:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_LP%A_84_29# 1 2 9 12 13 15 16 20 22 24 27 29 30
+ 34 35 37 38 39 40 41 44 48 50
r96 46 48 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.065 $Y=0.855
+ $X2=2.065 $Y2=0.485
r97 42 44 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.935 $Y=2.545
+ $X2=1.935 $Y2=2.845
r98 40 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.9 $Y=0.94
+ $X2=2.065 $Y2=0.855
r99 40 41 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=1.9 $Y=0.94
+ $X2=0.855 $Y2=0.94
r100 38 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.77 $Y=2.46
+ $X2=1.935 $Y2=2.545
r101 38 39 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.77 $Y=2.46
+ $X2=0.83 $Y2=2.46
r102 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.745 $Y=2.375
+ $X2=0.83 $Y2=2.46
r103 37 50 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.745 $Y=2.375
+ $X2=0.745 $Y2=1.555
r104 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.05 $X2=0.69 $Y2=1.05
r105 32 50 7.81933 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.39
+ $X2=0.69 $Y2=1.555
r106 32 34 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.69 $Y=1.39
+ $X2=0.69 $Y2=1.05
r107 31 41 16.4861 $w=1.17e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.855 $Y2=0.94
r108 31 34 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.69 $Y=1.025
+ $X2=0.69 $Y2=1.05
r109 28 35 36.8212 $w=4.35e-07 $l=2.88e-07 $layer=POLY_cond $X=0.637 $Y=1.338
+ $X2=0.637 $Y2=1.05
r110 28 29 47.0786 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.637 $Y=1.338
+ $X2=0.637 $Y2=1.555
r111 27 35 1.91777 $w=4.35e-07 $l=1.5e-08 $layer=POLY_cond $X=0.637 $Y=1.035
+ $X2=0.637 $Y2=1.05
r112 22 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.9 $Y=2.525
+ $X2=0.9 $Y2=2.845
r113 17 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=2.45
+ $X2=0.54 $Y2=2.45
r114 16 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.825 $Y=2.45
+ $X2=0.9 $Y2=2.525
r115 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.825 $Y=2.45
+ $X2=0.615 $Y2=2.45
r116 13 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.54 $Y=2.525
+ $X2=0.54 $Y2=2.45
r117 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=2.525
+ $X2=0.54 $Y2=2.845
r118 12 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.54 $Y=2.375
+ $X2=0.54 $Y2=2.45
r119 12 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.54 $Y=2.375
+ $X2=0.54 $Y2=1.555
r120 7 27 24.5823 $w=4.35e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=0.885
+ $X2=0.675 $Y2=1.035
r121 7 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.855 $Y=0.885
+ $X2=0.855 $Y2=0.485
r122 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.885
+ $X2=0.495 $Y2=0.485
r123 2 44 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=2.635 $X2=1.935 $Y2=2.845
r124 1 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.275 $X2=2.065 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP%A_200_367# 1 2 11 15 19 21 25 28 30 31 35 37
+ 41
c82 21 0 1.90523e-19 $X=3.845 $Y=2.12
r83 37 39 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.02 $Y=0.485
+ $X2=4.02 $Y2=0.715
r84 31 42 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=1.202 $Y=2 $X2=1.202
+ $Y2=2.165
r85 31 41 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=1.202 $Y=2 $X2=1.202
+ $Y2=1.835
r86 30 33 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.165 $Y=2 $X2=1.165
+ $Y2=2.12
r87 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165 $Y=2
+ $X2=1.165 $Y2=2
r88 28 35 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.1 $Y=2.035
+ $X2=4.015 $Y2=2.12
r89 28 39 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=4.1 $Y=2.035
+ $X2=4.1 $Y2=0.715
r90 23 35 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=2.205
+ $X2=4.015 $Y2=2.12
r91 23 25 21.693 $w=3.38e-07 $l=6.4e-07 $layer=LI1_cond $X=4.015 $Y=2.205
+ $X2=4.015 $Y2=2.845
r92 22 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=2.12
+ $X2=1.165 $Y2=2.12
r93 21 35 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.845 $Y=2.12
+ $X2=4.015 $Y2=2.12
r94 21 22 164.08 $w=1.68e-07 $l=2.515e-06 $layer=LI1_cond $X=3.845 $Y=2.12
+ $X2=1.33 $Y2=2.12
r95 17 19 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.215 $Y=0.95
+ $X2=1.46 $Y2=0.95
r96 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.46 $Y=0.875
+ $X2=1.46 $Y2=0.95
r97 13 15 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.46 $Y=0.875
+ $X2=1.46 $Y2=0.485
r98 11 42 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.33 $Y=2.845
+ $X2=1.33 $Y2=2.165
r99 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.215 $Y=1.025
+ $X2=1.215 $Y2=0.95
r100 7 41 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.215 $Y=1.025
+ $X2=1.215 $Y2=1.835
r101 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=2.635 $X2=4.01 $Y2=2.845
r102 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.88
+ $Y=0.275 $X2=4.02 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP%A1 3 7 9 10 13 14 18 21 22
c63 10 0 1.82988e-19 $X=1.83 $Y=1.28
r64 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.43
+ $X2=1.665 $Y2=1.595
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.43 $X2=1.665 $Y2=1.43
r66 18 22 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=1.665 $Y2=1.43
r67 14 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.565 $Y=1.13
+ $X2=2.565 $Y2=0.965
r68 13 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.565 $Y=1.13
+ $X2=2.565 $Y2=1.28
r69 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.565
+ $Y=1.13 $X2=2.565 $Y2=1.13
r70 11 22 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.665 $Y=1.365
+ $X2=1.665 $Y2=1.43
r71 10 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.83 $Y=1.28
+ $X2=1.665 $Y2=1.365
r72 9 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=1.28 $X2=2.565
+ $Y2=1.28
r73 9 10 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.4 $Y=1.28 $X2=1.83
+ $Y2=1.28
r74 7 26 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.505 $Y=0.485
+ $X2=2.505 $Y2=0.965
r75 3 24 640.957 $w=1.5e-07 $l=1.25e-06 $layer=POLY_cond $X=1.72 $Y=2.845
+ $X2=1.72 $Y2=1.595
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP%A0 1 3 8 12 14 15 16 21 23
c52 16 0 3.29388e-20 $X=3.12 $Y=1.665
c53 12 0 1.82988e-19 $X=2.115 $Y=0.88
r54 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.7
+ $X2=2.205 $Y2=1.865
r55 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.7
+ $X2=2.205 $Y2=1.535
r56 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.7 $X2=3.12
+ $Y2=1.7
r57 14 15 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.7 $X2=2.64
+ $Y2=1.7
r58 14 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.205
+ $Y=1.7 $X2=2.205 $Y2=1.7
r59 10 12 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.85 $Y=0.88
+ $X2=2.115 $Y2=0.88
r60 8 24 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.15 $Y=2.845
+ $X2=2.15 $Y2=1.865
r61 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.115 $Y=0.955
+ $X2=2.115 $Y2=0.88
r62 4 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.115 $Y=0.955
+ $X2=2.115 $Y2=1.535
r63 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=0.805
+ $X2=1.85 $Y2=0.88
r64 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.85 $Y=0.805 $X2=1.85
+ $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP%S 3 5 6 9 12 13 17 21 25 29 31 34 36 38 39
+ 43
c68 31 0 1.90523e-19 $X=3.03 $Y=1.79
c69 5 0 3.29388e-20 $X=2.97 $Y=2.18
r70 38 39 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.665
r71 38 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.36 $X2=3.57 $Y2=1.36
r72 35 43 37.2422 $w=5.1e-07 $l=3.55e-07 $layer=POLY_cond $X=3.615 $Y=1.715
+ $X2=3.615 $Y2=1.36
r73 35 36 7.86808 $w=5.1e-07 $l=7.5e-08 $layer=POLY_cond $X=3.615 $Y=1.715
+ $X2=3.615 $Y2=1.79
r74 34 43 1.57362 $w=5.1e-07 $l=1.5e-08 $layer=POLY_cond $X=3.615 $Y=1.345
+ $X2=3.615 $Y2=1.36
r75 19 34 24.7327 $w=5.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.62 $Y=1.195
+ $X2=3.62 $Y2=1.345
r76 19 29 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.805 $Y=1.195
+ $X2=3.805 $Y2=0.485
r77 19 21 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.445 $Y=1.195
+ $X2=3.445 $Y2=0.485
r78 15 36 37.3844 $w=5.1e-07 $l=7.5e-08 $layer=POLY_cond $X=3.615 $Y=1.865
+ $X2=3.615 $Y2=1.79
r79 15 25 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.795 $Y=1.865
+ $X2=3.795 $Y2=2.845
r80 15 17 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.435 $Y=1.865
+ $X2=3.435 $Y2=2.845
r81 14 31 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.12 $Y=1.79 $X2=3.03
+ $Y2=1.79
r82 13 36 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=3.36 $Y=1.79
+ $X2=3.615 $Y2=1.79
r83 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.36 $Y=1.79
+ $X2=3.12 $Y2=1.79
r84 11 31 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.045 $Y=1.865
+ $X2=3.03 $Y2=1.79
r85 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.045 $Y=1.865
+ $X2=3.045 $Y2=2.105
r86 7 31 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.015 $Y=1.715
+ $X2=3.03 $Y2=1.79
r87 7 9 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=3.015 $Y=1.715
+ $X2=3.015 $Y2=0.485
r88 5 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.97 $Y=2.18
+ $X2=3.045 $Y2=2.105
r89 5 6 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=2.97 $Y=2.18
+ $X2=2.615 $Y2=2.18
r90 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.54 $Y=2.255
+ $X2=2.615 $Y2=2.18
r91 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.54 $Y=2.255 $X2=2.54
+ $Y2=2.845
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP%X 1 2 9 12 13 14 15 16 17
r20 16 17 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=2.035
+ $X2=0.235 $Y2=2.405
r21 15 16 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=2.035
r22 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r23 13 14 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=1.295
r24 13 39 10.0839 $w=2.38e-07 $l=2.1e-07 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=0.715
r25 12 39 8.90991 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.28 $Y=0.485
+ $X2=0.28 $Y2=0.715
r26 10 17 10.0839 $w=2.38e-07 $l=2.1e-07 $layer=LI1_cond $X=0.235 $Y=2.615
+ $X2=0.235 $Y2=2.405
r27 9 10 8.55704 $w=3.73e-07 $l=2.3e-07 $layer=LI1_cond $X=0.302 $Y=2.845
+ $X2=0.302 $Y2=2.615
r28 2 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=2.635 $X2=0.325 $Y2=2.845
r29 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.275 $X2=0.28 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP%VPWR 1 2 9 11 15 17 19 29 30 33 36
r46 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=4.08
+ $Y2=3.33
r52 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=3.33
+ $X2=2.755 $Y2=3.33
r54 24 26 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.92 $Y=3.33 $X2=3.12
+ $Y2=3.33
r55 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=1.115 $Y2=3.33
r58 19 21 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 17 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=3.245
+ $X2=2.755 $Y2=3.33
r62 13 15 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.755 $Y=3.245
+ $X2=2.755 $Y2=2.845
r63 12 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=3.33
+ $X2=1.115 $Y2=3.33
r64 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=2.755 $Y2=3.33
r65 11 12 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=1.28 $Y2=3.33
r66 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=3.245
+ $X2=1.115 $Y2=3.33
r67 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.115 $Y=3.245
+ $X2=1.115 $Y2=2.895
r68 2 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=2.635 $X2=2.755 $Y2=2.845
r69 1 9 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=2.635 $X2=1.115 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_LP%VGND 1 2 9 11 15 17 19 26 27 30 33
r45 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r48 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r49 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.23
+ $Y2=0
r50 24 26 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=4.08
+ $Y2=0
r51 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r52 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r54 19 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r55 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r56 17 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r57 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=0.085
+ $X2=3.23 $Y2=0
r58 13 15 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.23 $Y=0.085 $X2=3.23
+ $Y2=0.485
r59 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r60 11 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=3.23
+ $Y2=0
r61 11 12 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=3.065 $Y=0 $X2=1.235
+ $Y2=0
r62 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r63 7 9 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.47
r64 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.275 $X2=3.23 $Y2=0.485
r65 1 9 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.275 $X2=1.07 $Y2=0.47
.ends

