* File: sky130_fd_sc_lp__sdfrtn_1.spice
* Created: Wed Sep  2 10:34:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrtn_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfrtn_1  VNB VPB SCD SCE D RESET_B CLK_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK_N	CLK_N
* RESET_B	RESET_B
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1039 N_A_113_63#_M1039_d N_SCE_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 noxref_25 N_SCD_M1026_g N_noxref_24_M1026_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1028 N_A_229_491#_M1028_d N_SCE_M1028_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.12305 AS=0.0441 PD=1.04 PS=0.63 NRD=34.284 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 noxref_26 N_D_M1010_g N_A_229_491#_M1028_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.12305 PD=0.69 PS=1.04 NRD=22.848 NRS=34.284 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 N_noxref_24_M1015_d N_A_113_63#_M1015_g noxref_26 VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0567 PD=0.81 PS=0.69 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.6 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_RESET_B_M1034_g N_noxref_24_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.122292 AS=0.0819 PD=0.95 PS=0.81 NRD=34.284 NRS=31.428 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1023 N_A_857_367#_M1023_d N_CLK_N_M1023_g N_VGND_M1034_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.244583 PD=2.25 PS=1.9 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75001.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1019 N_A_1080_47#_M1019_d N_A_857_367#_M1019_g N_VGND_M1019_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.3679 AS=0.2394 PD=2.7 PS=2.25 NRD=17.136 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1020 N_A_1278_529#_M1020_d N_A_1080_47#_M1020_g N_A_229_491#_M1020_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.2247 PD=0.7 PS=1.91 NRD=0 NRS=74.28 M=1
+ R=2.8 SA=75000.5 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1008 A_1437_127# N_A_857_367#_M1008_g N_A_1278_529#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75004.5 A=0.063 P=1.14 MULT=1
MM1007 A_1509_127# N_A_1406_399#_M1007_g A_1437_127# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75004.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_1509_127# VNB NSHORT L=0.15 W=0.42
+ AD=0.175588 AS=0.0441 PD=1.25208 PS=0.63 NRD=103.728 NRS=14.28 M=1 R=2.8
+ SA=75001.6 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_1406_399#_M1001_d N_A_1278_529#_M1001_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.163925 AS=0.267562 PD=1.155 PS=1.90792 NRD=21.552
+ NRS=68.064 M=1 R=4.26667 SA=75001.7 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1016 N_A_1870_127#_M1016_d N_A_857_367#_M1016_g N_A_1406_399#_M1001_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.221102 AS=0.163925 PD=1.50943 PS=1.155 NRD=40.308
+ NRS=21.552 M=1 R=4.26667 SA=75002.3 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1017 A_2022_127# N_A_1080_47#_M1017_g N_A_1870_127#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.145098 PD=0.63 PS=0.990566 NRD=14.28 NRS=33.564 M=1
+ R=2.8 SA=75003.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_2064_101#_M1029_g A_2022_127# VNB NSHORT L=0.15 W=0.42
+ AD=0.1071 AS=0.0441 PD=0.93 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8 SA=75004.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 A_2226_127# N_RESET_B_M1002_g N_VGND_M1029_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1071 PD=0.63 PS=0.93 NRD=14.28 NRS=32.856 M=1 R=2.8 SA=75004.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_2064_101#_M1030_d N_A_1870_127#_M1030_g A_2226_127# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75005.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_1870_127#_M1011_g N_A_2370_351#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=9.996 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1031 N_Q_M1031_d N_A_2370_351#_M1031_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=4.284 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_A_113_63#_M1021_d N_SCE_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1032 A_312_491# N_A_113_63#_M1032_g N_A_229_491#_M1032_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1037 N_VPWR_M1037_d N_SCD_M1037_g A_312_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2663 AS=0.0672 PD=1.48 PS=0.85 NRD=19.9955 NRS=15.3857 M=1 R=4.26667
+ SA=75000.6 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1014 A_562_491# N_SCE_M1014_g N_VPWR_M1037_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.2663 PD=0.85 PS=1.48 NRD=15.3857 NRS=19.9955 M=1 R=4.26667
+ SA=75001.4 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1018 N_A_229_491#_M1018_d N_D_M1018_g A_562_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=15.3857 NRS=15.3857 M=1 R=4.26667
+ SA=75001.8 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_RESET_B_M1000_g N_A_229_491#_M1018_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.146964 AS=0.1248 PD=1.13516 PS=1.03 NRD=21.5321 NRS=18.4589 M=1
+ R=4.26667 SA=75002.3 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1035 N_A_857_367#_M1035_d N_CLK_N_M1035_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.289336 PD=3.05 PS=2.23484 NRD=0 NRS=11.7215 M=1 R=8.4
+ SA=75001.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1022 N_A_1080_47#_M1022_d N_A_857_367#_M1022_g N_VPWR_M1022_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_1278_529#_M1005_d N_A_857_367#_M1005_g N_A_229_491#_M1005_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1027 A_1364_529# N_A_1080_47#_M1027_g N_A_1278_529#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_A_1406_399#_M1036_g A_1364_529# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_1278_529#_M1003_d N_RESET_B_M1003_g N_VPWR_M1036_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 N_A_1406_399#_M1038_d N_A_1278_529#_M1038_g N_VPWR_M1038_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.3679 PD=1.12 PS=2.7 NRD=0 NRS=28.1316 M=1 R=5.6
+ SA=75000.3 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1006 N_A_1870_127#_M1006_d N_A_1080_47#_M1006_g N_A_1406_399#_M1038_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1792 AS=0.1176 PD=1.62 PS=1.12 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.8 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1024 A_2022_533# N_A_857_367#_M1024_g N_A_1870_127#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=74.2493 M=1 R=2.8
+ SA=75001.3 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_2064_101#_M1012_g A_2022_533# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.10185 AS=0.0441 PD=0.905 PS=0.63 NRD=44.5417 NRS=23.443 M=1 R=2.8
+ SA=75001.6 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1033 N_A_2064_101#_M1033_d N_RESET_B_M1033_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.10185 PD=0.7 PS=0.905 NRD=0 NRS=51.5943 M=1 R=2.8
+ SA=75002.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_1870_127#_M1013_g N_A_2064_101#_M1033_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_1870_127#_M1004_g N_A_2370_351#_M1004_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.174989 AS=0.1696 PD=1.21937 PS=1.81 NRD=40.779 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1025 N_Q_M1025_d N_A_2370_351#_M1025_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.344511 PD=3.09 PS=2.40063 NRD=3.1126 NRS=9.3772 M=1
+ R=8.4 SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.8651 P=31.53
*
.include "sky130_fd_sc_lp__sdfrtn_1.pxi.spice"
*
.ends
*
*
