# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.590000 1.210000 2.075000 2.145000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.235000 0.375000 9.505000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.255000 0.355000 8.545000 2.205000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.425000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.670000 ;
        RECT 1.755000  0.085000 2.075000 0.975000 ;
        RECT 3.610000  0.085000 4.335000 0.915000 ;
        RECT 6.050000  0.085000 6.380000 0.955000 ;
        RECT 7.775000  0.085000 8.085000 1.230000 ;
        RECT 8.745000  0.085000 9.015000 1.255000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.600000 3.415000 ;
        RECT 0.095000 2.320000 0.390000 3.245000 ;
        RECT 1.495000 2.655000 1.735000 3.245000 ;
        RECT 3.945000 2.765000 4.275000 3.245000 ;
        RECT 6.080000 1.975000 6.410000 3.245000 ;
        RECT 7.785000 2.715000 8.115000 3.245000 ;
        RECT 8.805000 2.785000 9.015000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.560000 2.320000 0.795000 2.990000 ;
      RECT 0.595000 0.450000 0.875000 1.215000 ;
      RECT 0.595000 1.215000 1.040000 1.885000 ;
      RECT 0.595000 1.885000 0.795000 2.320000 ;
      RECT 1.045000 2.295000 1.420000 2.315000 ;
      RECT 1.045000 2.315000 2.075000 2.485000 ;
      RECT 1.045000 2.485000 1.325000 2.965000 ;
      RECT 1.210000 0.640000 1.420000 2.295000 ;
      RECT 1.905000 2.485000 2.075000 2.865000 ;
      RECT 1.905000 2.865000 3.300000 3.075000 ;
      RECT 2.245000 0.635000 2.695000 0.965000 ;
      RECT 2.245000 0.965000 2.435000 2.695000 ;
      RECT 2.605000 1.555000 4.460000 1.725000 ;
      RECT 2.605000 1.725000 2.775000 2.365000 ;
      RECT 2.605000 2.365000 2.960000 2.695000 ;
      RECT 2.865000 0.635000 3.160000 1.555000 ;
      RECT 2.945000 1.895000 3.300000 2.155000 ;
      RECT 3.130000 2.155000 3.300000 2.415000 ;
      RECT 3.130000 2.415000 5.035000 2.585000 ;
      RECT 3.130000 2.585000 3.300000 2.865000 ;
      RECT 3.495000 1.895000 4.695000 2.235000 ;
      RECT 3.545000 1.085000 4.695000 1.255000 ;
      RECT 3.545000 1.255000 3.875000 1.385000 ;
      RECT 4.130000 1.425000 4.460000 1.555000 ;
      RECT 4.505000 0.585000 4.695000 1.085000 ;
      RECT 4.865000 1.225000 5.095000 1.555000 ;
      RECT 4.865000 1.555000 5.035000 2.415000 ;
      RECT 5.010000 0.640000 5.435000 0.995000 ;
      RECT 5.205000 1.875000 5.465000 2.750000 ;
      RECT 5.265000 0.995000 5.435000 1.125000 ;
      RECT 5.265000 1.125000 6.685000 1.295000 ;
      RECT 5.265000 1.295000 5.465000 1.875000 ;
      RECT 5.895000 1.485000 6.225000 1.635000 ;
      RECT 5.895000 1.635000 7.265000 1.650000 ;
      RECT 5.895000 1.650000 7.035000 1.805000 ;
      RECT 6.435000 1.295000 6.685000 1.455000 ;
      RECT 6.550000 0.355000 6.890000 0.775000 ;
      RECT 6.550000 0.775000 7.035000 0.955000 ;
      RECT 6.580000 1.805000 7.035000 2.375000 ;
      RECT 6.580000 2.375000 9.050000 2.545000 ;
      RECT 6.580000 2.545000 6.875000 2.755000 ;
      RECT 6.865000 0.955000 7.035000 1.320000 ;
      RECT 6.865000 1.320000 7.265000 1.635000 ;
      RECT 7.060000 0.265000 7.385000 0.595000 ;
      RECT 7.215000 0.595000 7.385000 0.830000 ;
      RECT 7.215000 0.830000 7.605000 1.040000 ;
      RECT 7.260000 1.875000 7.605000 2.205000 ;
      RECT 7.435000 1.040000 7.605000 1.875000 ;
      RECT 8.720000 1.425000 9.050000 2.375000 ;
  END
END sky130_fd_sc_lp__dfxbp_1
