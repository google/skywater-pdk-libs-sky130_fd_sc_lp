* File: sky130_fd_sc_lp__or2_0.spice
* Created: Wed Sep  2 10:28:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2_0.pex.spice"
.subckt sky130_fd_sc_lp__or2_0  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1002 N_A_76_473#_M1002_d N_B_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_76_473#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_76_473#_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 A_159_473# N_B_M1000_g N_A_76_473#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_159_473# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.143711 AS=0.0504 PD=0.998491 PS=0.66 NRD=56.2829 NRS=30.4759 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_76_473#_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.218989 PD=1.81 PS=1.52151 NRD=0 NRS=16.154 M=1 R=4.26667
+ SA=75001 SB=75000.2 A=0.096 P=1.58 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_50 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__or2_0.pxi.spice"
*
.ends
*
*
