* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1237_55# a_794_47# a_1327_415# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1327_415# a_1365_29# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_1365_29# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_208_481# D a_244_121# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_1888_463# a_963_47# a_1998_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 Q a_2686_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VPWR a_794_47# a_963_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VPWR a_2686_131# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND SCD a_172_121# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_1998_463# a_2214_99# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR a_1237_55# a_1365_29# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_1998_463# a_794_47# a_1781_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 Q a_2686_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_244_121# D a_330_121# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_244_121# a_794_47# a_1237_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_2159_125# a_2214_99# a_2244_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1365_29# a_1237_55# a_1608_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR SCE a_358_429# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_2686_131# a_1998_463# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_244_121# a_963_47# a_1237_55# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_1323_55# a_1365_29# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VGND a_1237_55# a_1933_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_330_121# a_358_429# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_794_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VGND a_794_47# a_963_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_2686_131# a_1998_463# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_244_121# a_358_429# a_39_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 VPWR SET_B a_1998_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_2244_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1888_463# a_2214_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VPWR SCE a_208_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_1608_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_794_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 VPWR a_1237_55# a_1781_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X34 a_1933_125# a_963_47# a_1998_463# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 VGND SCE a_358_429# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_1237_55# a_963_47# a_1323_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VGND a_2686_131# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 a_39_481# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 a_172_121# SCE a_244_121# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_1998_463# a_794_47# a_2159_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 VGND a_1998_463# a_2214_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
