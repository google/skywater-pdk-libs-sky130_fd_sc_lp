* File: sky130_fd_sc_lp__iso1n_lp2.pxi.spice
* Created: Fri Aug 28 10:41:05 2020
* 
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%SLEEP_B N_SLEEP_B_c_63_n N_SLEEP_B_M1001_g
+ N_SLEEP_B_c_64_n N_SLEEP_B_c_65_n N_SLEEP_B_M1000_g N_SLEEP_B_c_66_n
+ N_SLEEP_B_M1006_g N_SLEEP_B_c_67_n SLEEP_B N_SLEEP_B_c_68_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP2%SLEEP_B
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%A_27_109# N_A_27_109#_M1001_s
+ N_A_27_109#_M1000_s N_A_27_109#_M1008_g N_A_27_109#_M1007_g
+ N_A_27_109#_M1004_g N_A_27_109#_c_108_n N_A_27_109#_c_116_n
+ N_A_27_109#_c_109_n N_A_27_109#_c_117_n N_A_27_109#_c_110_n
+ N_A_27_109#_c_111_n N_A_27_109#_c_118_n N_A_27_109#_c_112_n
+ N_A_27_109#_c_113_n N_A_27_109#_c_114_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP2%A_27_109#
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%A N_A_M1002_g N_A_M1011_g N_A_M1009_g A A
+ N_A_c_188_n PM_SKY130_FD_SC_LP__ISO1N_LP2%A
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%A_350_109# N_A_350_109#_M1004_d
+ N_A_350_109#_M1002_d N_A_350_109#_M1010_g N_A_350_109#_M1003_g
+ N_A_350_109#_M1005_g N_A_350_109#_c_228_n N_A_350_109#_c_233_n
+ N_A_350_109#_c_234_n N_A_350_109#_c_229_n N_A_350_109#_c_230_n
+ N_A_350_109#_c_231_n N_A_350_109#_c_236_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP2%A_350_109#
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%VPWR N_VPWR_M1000_d N_VPWR_M1003_s
+ N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_299_n VPWR
+ N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_295_n N_VPWR_c_303_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP2%VPWR
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%X N_X_M1005_d N_X_M1003_d X X X X X N_X_c_330_n
+ X X PM_SKY130_FD_SC_LP__ISO1N_LP2%X
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%KAGND N_KAGND_M1006_d N_KAGND_M1009_d KAGND
+ N_KAGND_c_349_n N_KAGND_c_350_n N_KAGND_c_351_n N_KAGND_c_352_n
+ PM_SKY130_FD_SC_LP__ISO1N_LP2%KAGND
x_PM_SKY130_FD_SC_LP__ISO1N_LP2%VGND VGND N_VGND_c_400_n N_VGND_c_401_n VGND
+ PM_SKY130_FD_SC_LP__ISO1N_LP2%VGND
cc_1 VNB N_SLEEP_B_c_63_n 0.0168134f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.04
cc_2 VNB N_SLEEP_B_c_64_n 0.018582f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_3 VNB N_SLEEP_B_c_65_n 0.0148835f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.115
cc_4 VNB N_SLEEP_B_c_66_n 0.0127833f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.04
cc_5 VNB N_SLEEP_B_c_67_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.115
cc_6 VNB N_SLEEP_B_c_68_n 0.0204036f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.68
cc_7 VNB N_A_27_109#_M1008_g 0.0194021f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.545
cc_8 VNB N_A_27_109#_M1004_g 0.0195709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_109#_c_108_n 0.0298351f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.68
cc_10 VNB N_A_27_109#_c_109_n 0.023802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_109#_c_110_n 0.0128314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_109#_c_111_n 0.0132078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_109#_c_112_n 0.0150831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_109#_c_113_n 0.00140221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_109#_c_114_n 0.0301343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_M1011_g 0.0202362f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.115
cc_17 VNB N_A_M1009_g 0.0189609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A 0.00326145f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.755
cc_19 VNB N_A_c_188_n 0.0750523f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.68
cc_20 VNB N_A_350_109#_M1010_g 0.0194066f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.545
cc_21 VNB N_A_350_109#_M1005_g 0.0233516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_350_109#_c_228_n 0.00684374f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.68
cc_23 VNB N_A_350_109#_c_229_n 5.62227e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_350_109#_c_230_n 0.0487169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_350_109#_c_231_n 0.00316756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_295_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0347504f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.115
cc_28 VNB N_X_c_330_n 0.0172805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_KAGND_c_349_n 0.0169074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_KAGND_c_350_n 0.013451f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.68
cc_31 VNB N_KAGND_c_351_n 0.0214252f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.68
cc_32 VNB N_KAGND_c_352_n 0.0300475f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.68
cc_33 VNB N_VGND_c_400_n 0.227491f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_34 VNB N_VGND_c_401_n 0.101553f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.845
cc_35 VPB N_SLEEP_B_M1000_g 0.0339923f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.545
cc_36 VPB N_SLEEP_B_c_68_n 0.0265795f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.68
cc_37 VPB N_A_27_109#_M1007_g 0.0295722f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.755
cc_38 VPB N_A_27_109#_c_116_n 0.0139274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_109#_c_117_n 0.0429724f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_109#_c_118_n 0.0201745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_109#_c_112_n 0.0180068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_27_109#_c_113_n 0.001264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_27_109#_c_114_n 9.90415e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_M1002_g 0.0407024f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.755
cc_45 VPB N_A_c_188_n 0.0123468f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.68
cc_46 VPB N_A_350_109#_M1003_g 0.0392909f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.755
cc_47 VPB N_A_350_109#_c_233_n 0.0300703f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.68
cc_48 VPB N_A_350_109#_c_234_n 0.0315384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_350_109#_c_230_n 0.027476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_350_109#_c_236_n 0.00137249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_296_n 0.0146662f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.545
cc_52 VPB N_VPWR_c_297_n 0.0236277f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.115
cc_53 VPB N_VPWR_c_298_n 0.0459711f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.68
cc_54 VPB N_VPWR_c_299_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.68
cc_55 VPB N_VPWR_c_300_n 0.0255379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_301_n 0.0192431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_295_n 0.0890167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_303_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB X 0.0190114f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.115
cc_60 VPB X 0.035517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB X 0.00736113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 N_SLEEP_B_c_66_n N_A_27_109#_M1008_g 0.0178481f $X=0.855 $Y=1.04 $X2=0
+ $Y2=0
cc_63 N_SLEEP_B_c_68_n N_A_27_109#_M1007_g 0.0149412f $X=0.805 $Y=1.68 $X2=0
+ $Y2=0
cc_64 N_SLEEP_B_c_64_n N_A_27_109#_c_108_n 0.00271235f $X=0.495 $Y=1.515 $X2=0
+ $Y2=0
cc_65 N_SLEEP_B_c_65_n N_A_27_109#_c_108_n 0.0013897f $X=0.78 $Y=1.115 $X2=0
+ $Y2=0
cc_66 N_SLEEP_B_c_63_n N_A_27_109#_c_109_n 0.00911088f $X=0.495 $Y=1.04 $X2=0
+ $Y2=0
cc_67 N_SLEEP_B_c_66_n N_A_27_109#_c_109_n 8.53265e-19 $X=0.855 $Y=1.04 $X2=0
+ $Y2=0
cc_68 N_SLEEP_B_c_67_n N_A_27_109#_c_109_n 0.00834731f $X=0.495 $Y=1.115 $X2=0
+ $Y2=0
cc_69 N_SLEEP_B_c_64_n N_A_27_109#_c_110_n 0.00609799f $X=0.495 $Y=1.515 $X2=0
+ $Y2=0
cc_70 N_SLEEP_B_c_65_n N_A_27_109#_c_110_n 0.0104164f $X=0.78 $Y=1.115 $X2=0
+ $Y2=0
cc_71 N_SLEEP_B_c_67_n N_A_27_109#_c_110_n 0.00300872f $X=0.495 $Y=1.115 $X2=0
+ $Y2=0
cc_72 SLEEP_B N_A_27_109#_c_110_n 0.0235108f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_73 N_SLEEP_B_c_68_n N_A_27_109#_c_110_n 0.00405919f $X=0.805 $Y=1.68 $X2=0
+ $Y2=0
cc_74 N_SLEEP_B_c_64_n N_A_27_109#_c_111_n 0.00447049f $X=0.495 $Y=1.515 $X2=0
+ $Y2=0
cc_75 N_SLEEP_B_c_67_n N_A_27_109#_c_111_n 5.63939e-19 $X=0.495 $Y=1.115 $X2=0
+ $Y2=0
cc_76 N_SLEEP_B_M1000_g N_A_27_109#_c_118_n 0.00107346f $X=0.805 $Y=2.545 $X2=0
+ $Y2=0
cc_77 SLEEP_B N_A_27_109#_c_118_n 0.00961287f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_78 N_SLEEP_B_c_68_n N_A_27_109#_c_118_n 0.00708073f $X=0.805 $Y=1.68 $X2=0
+ $Y2=0
cc_79 N_SLEEP_B_c_64_n N_A_27_109#_c_112_n 0.0139429f $X=0.495 $Y=1.515 $X2=0
+ $Y2=0
cc_80 N_SLEEP_B_M1000_g N_A_27_109#_c_112_n 0.00370596f $X=0.805 $Y=2.545 $X2=0
+ $Y2=0
cc_81 SLEEP_B N_A_27_109#_c_112_n 0.0203945f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_82 N_SLEEP_B_c_64_n N_A_27_109#_c_113_n 4.46737e-19 $X=0.495 $Y=1.515 $X2=0
+ $Y2=0
cc_83 SLEEP_B N_A_27_109#_c_113_n 0.0139191f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_84 N_SLEEP_B_c_68_n N_A_27_109#_c_113_n 0.00135236f $X=0.805 $Y=1.68 $X2=0
+ $Y2=0
cc_85 SLEEP_B N_A_27_109#_c_114_n 0.00101513f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_86 N_SLEEP_B_c_68_n N_A_27_109#_c_114_n 0.0174467f $X=0.805 $Y=1.68 $X2=0
+ $Y2=0
cc_87 N_SLEEP_B_M1000_g N_VPWR_c_296_n 0.0226892f $X=0.805 $Y=2.545 $X2=0 $Y2=0
cc_88 N_SLEEP_B_M1000_g N_VPWR_c_300_n 0.00802402f $X=0.805 $Y=2.545 $X2=0 $Y2=0
cc_89 N_SLEEP_B_M1000_g N_VPWR_c_295_n 0.0150852f $X=0.805 $Y=2.545 $X2=0 $Y2=0
cc_90 N_SLEEP_B_c_63_n N_KAGND_c_349_n 0.00358937f $X=0.495 $Y=1.04 $X2=0 $Y2=0
cc_91 N_SLEEP_B_c_66_n N_KAGND_c_349_n 0.0159665f $X=0.855 $Y=1.04 $X2=0 $Y2=0
cc_92 N_SLEEP_B_c_63_n N_KAGND_c_352_n 0.00463047f $X=0.495 $Y=1.04 $X2=0 $Y2=0
cc_93 N_SLEEP_B_c_65_n N_KAGND_c_352_n 6.11331e-19 $X=0.78 $Y=1.115 $X2=0 $Y2=0
cc_94 N_SLEEP_B_c_63_n N_VGND_c_400_n 0.00293597f $X=0.495 $Y=1.04 $X2=0 $Y2=0
cc_95 N_SLEEP_B_c_63_n N_VGND_c_401_n 0.00441768f $X=0.495 $Y=1.04 $X2=0 $Y2=0
cc_96 N_SLEEP_B_c_66_n N_VGND_c_401_n 6.46133e-19 $X=0.855 $Y=1.04 $X2=0 $Y2=0
cc_97 N_A_27_109#_c_116_n N_A_M1002_g 0.0425499f $X=1.335 $Y=1.835 $X2=0 $Y2=0
cc_98 N_A_27_109#_M1004_g N_A_M1011_g 0.0176841f $X=1.675 $Y=0.755 $X2=0 $Y2=0
cc_99 N_A_27_109#_c_108_n N_A_c_188_n 0.0076954f $X=1.675 $Y=1.24 $X2=0 $Y2=0
cc_100 N_A_27_109#_c_113_n N_A_c_188_n 3.2833e-19 $X=1.335 $Y=1.33 $X2=0 $Y2=0
cc_101 N_A_27_109#_c_114_n N_A_c_188_n 0.0465204f $X=1.335 $Y=1.33 $X2=0 $Y2=0
cc_102 N_A_27_109#_M1008_g N_A_350_109#_c_228_n 9.51545e-19 $X=1.285 $Y=0.755
+ $X2=0 $Y2=0
cc_103 N_A_27_109#_M1004_g N_A_350_109#_c_228_n 0.00502952f $X=1.675 $Y=0.755
+ $X2=0 $Y2=0
cc_104 N_A_27_109#_c_108_n N_A_350_109#_c_228_n 0.00510417f $X=1.675 $Y=1.24
+ $X2=0 $Y2=0
cc_105 N_A_27_109#_c_113_n N_A_350_109#_c_228_n 0.0345812f $X=1.335 $Y=1.33
+ $X2=0 $Y2=0
cc_106 N_A_27_109#_c_114_n N_A_350_109#_c_228_n 0.00269832f $X=1.335 $Y=1.33
+ $X2=0 $Y2=0
cc_107 N_A_27_109#_M1007_g N_A_350_109#_c_233_n 0.00808597f $X=1.375 $Y=2.545
+ $X2=0 $Y2=0
cc_108 N_A_27_109#_M1008_g N_A_350_109#_c_231_n 4.37216e-19 $X=1.285 $Y=0.755
+ $X2=0 $Y2=0
cc_109 N_A_27_109#_M1004_g N_A_350_109#_c_231_n 0.00619682f $X=1.675 $Y=0.755
+ $X2=0 $Y2=0
cc_110 N_A_27_109#_c_116_n N_A_350_109#_c_236_n 0.0013215f $X=1.335 $Y=1.835
+ $X2=0 $Y2=0
cc_111 N_A_27_109#_c_113_n N_A_350_109#_c_236_n 0.0121722f $X=1.335 $Y=1.33
+ $X2=0 $Y2=0
cc_112 N_A_27_109#_M1007_g N_VPWR_c_296_n 0.00332866f $X=1.375 $Y=2.545 $X2=0
+ $Y2=0
cc_113 N_A_27_109#_c_116_n N_VPWR_c_296_n 4.86308e-19 $X=1.335 $Y=1.835 $X2=0
+ $Y2=0
cc_114 N_A_27_109#_c_118_n N_VPWR_c_296_n 0.0273824f $X=0.54 $Y=2.19 $X2=0 $Y2=0
cc_115 N_A_27_109#_c_113_n N_VPWR_c_296_n 0.00515663f $X=1.335 $Y=1.33 $X2=0
+ $Y2=0
cc_116 N_A_27_109#_M1007_g N_VPWR_c_298_n 0.00893366f $X=1.375 $Y=2.545 $X2=0
+ $Y2=0
cc_117 N_A_27_109#_c_117_n N_VPWR_c_300_n 0.0342516f $X=0.54 $Y=2.9 $X2=0 $Y2=0
cc_118 N_A_27_109#_M1007_g N_VPWR_c_295_n 0.0164524f $X=1.375 $Y=2.545 $X2=0
+ $Y2=0
cc_119 N_A_27_109#_c_117_n N_VPWR_c_295_n 0.0196561f $X=0.54 $Y=2.9 $X2=0 $Y2=0
cc_120 N_A_27_109#_M1008_g N_KAGND_c_349_n 0.0166532f $X=1.285 $Y=0.755 $X2=0
+ $Y2=0
cc_121 N_A_27_109#_M1004_g N_KAGND_c_349_n 0.00368399f $X=1.675 $Y=0.755 $X2=0
+ $Y2=0
cc_122 N_A_27_109#_c_108_n N_KAGND_c_349_n 3.10624e-19 $X=1.675 $Y=1.24 $X2=0
+ $Y2=0
cc_123 N_A_27_109#_c_109_n N_KAGND_c_349_n 0.0118897f $X=0.28 $Y=0.755 $X2=0
+ $Y2=0
cc_124 N_A_27_109#_c_110_n N_KAGND_c_349_n 0.0310664f $X=1.17 $Y=1.25 $X2=0
+ $Y2=0
cc_125 N_A_27_109#_c_113_n N_KAGND_c_349_n 0.016937f $X=1.335 $Y=1.33 $X2=0
+ $Y2=0
cc_126 N_A_27_109#_M1004_g N_KAGND_c_350_n 0.00541012f $X=1.675 $Y=0.755 $X2=0
+ $Y2=0
cc_127 N_A_27_109#_M1004_g N_KAGND_c_352_n 0.00746866f $X=1.675 $Y=0.755 $X2=0
+ $Y2=0
cc_128 N_A_27_109#_c_109_n N_KAGND_c_352_n 0.0323241f $X=0.28 $Y=0.755 $X2=0
+ $Y2=0
cc_129 N_A_27_109#_c_110_n N_KAGND_c_352_n 0.0108315f $X=1.17 $Y=1.25 $X2=0
+ $Y2=0
cc_130 N_A_27_109#_c_113_n N_KAGND_c_352_n 0.00502324f $X=1.335 $Y=1.33 $X2=0
+ $Y2=0
cc_131 N_A_27_109#_c_109_n N_VGND_c_400_n 0.00142664f $X=0.28 $Y=0.755 $X2=0
+ $Y2=0
cc_132 N_A_27_109#_M1008_g N_VGND_c_401_n 6.46133e-19 $X=1.285 $Y=0.755 $X2=0
+ $Y2=0
cc_133 N_A_27_109#_M1004_g N_VGND_c_401_n 6.46133e-19 $X=1.675 $Y=0.755 $X2=0
+ $Y2=0
cc_134 N_A_27_109#_c_109_n N_VGND_c_401_n 0.00876524f $X=0.28 $Y=0.755 $X2=0
+ $Y2=0
cc_135 N_A_M1009_g N_A_350_109#_M1010_g 0.017228f $X=2.545 $Y=0.755 $X2=0 $Y2=0
cc_136 A N_A_350_109#_M1010_g 0.00246135f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A_c_188_n N_A_350_109#_M1010_g 0.0212527f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_138 N_A_M1011_g N_A_350_109#_c_228_n 0.00352672f $X=2.185 $Y=0.755 $X2=0
+ $Y2=0
cc_139 A N_A_350_109#_c_228_n 0.0251831f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A_c_188_n N_A_350_109#_c_228_n 0.0138392f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_141 N_A_M1002_g N_A_350_109#_c_233_n 0.0390928f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_142 A N_A_350_109#_c_234_n 0.0333494f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A_c_188_n N_A_350_109#_c_234_n 0.00994677f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_144 A N_A_350_109#_c_229_n 0.0258605f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A_c_188_n N_A_350_109#_c_229_n 0.00128478f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_146 N_A_c_188_n N_A_350_109#_c_230_n 0.00444435f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_147 N_A_M1011_g N_A_350_109#_c_231_n 0.0021581f $X=2.185 $Y=0.755 $X2=0 $Y2=0
cc_148 A N_A_350_109#_c_231_n 7.35267e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A_c_188_n N_A_350_109#_c_231_n 0.00602809f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_150 N_A_M1002_g N_A_350_109#_c_236_n 0.00714529f $X=1.865 $Y=2.545 $X2=0
+ $Y2=0
cc_151 A N_A_350_109#_c_236_n 0.0192162f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A_c_188_n N_A_350_109#_c_236_n 0.0212357f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_VPWR_c_298_n 0.00545907f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_VPWR_c_295_n 0.00825001f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_155 N_A_M1011_g N_KAGND_c_350_n 0.00545157f $X=2.185 $Y=0.755 $X2=0 $Y2=0
cc_156 N_A_M1011_g N_KAGND_c_351_n 0.00377907f $X=2.185 $Y=0.755 $X2=0 $Y2=0
cc_157 N_A_M1009_g N_KAGND_c_351_n 0.0162067f $X=2.545 $Y=0.755 $X2=0 $Y2=0
cc_158 A N_KAGND_c_351_n 0.0236868f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A_c_188_n N_KAGND_c_351_n 0.0016217f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_160 N_A_M1011_g N_KAGND_c_352_n 0.00652703f $X=2.185 $Y=0.755 $X2=0 $Y2=0
cc_161 A N_KAGND_c_352_n 0.0137584f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A_c_188_n N_KAGND_c_352_n 0.00190945f $X=2.525 $Y=1.33 $X2=0 $Y2=0
cc_163 N_A_M1011_g N_VGND_c_401_n 6.46133e-19 $X=2.185 $Y=0.755 $X2=0 $Y2=0
cc_164 N_A_M1009_g N_VGND_c_401_n 6.46133e-19 $X=2.545 $Y=0.755 $X2=0 $Y2=0
cc_165 N_A_350_109#_c_233_n N_VPWR_c_296_n 0.00165396f $X=2.13 $Y=2.19 $X2=0
+ $Y2=0
cc_166 N_A_350_109#_M1003_g N_VPWR_c_297_n 0.0249766f $X=3.285 $Y=2.545 $X2=0
+ $Y2=0
cc_167 N_A_350_109#_c_233_n N_VPWR_c_297_n 0.0396681f $X=2.13 $Y=2.19 $X2=0
+ $Y2=0
cc_168 N_A_350_109#_c_234_n N_VPWR_c_297_n 0.0273651f $X=2.935 $Y=1.76 $X2=0
+ $Y2=0
cc_169 N_A_350_109#_c_230_n N_VPWR_c_297_n 0.00269508f $X=3.1 $Y=1.34 $X2=0
+ $Y2=0
cc_170 N_A_350_109#_c_233_n N_VPWR_c_298_n 0.0394541f $X=2.13 $Y=2.19 $X2=0
+ $Y2=0
cc_171 N_A_350_109#_M1003_g N_VPWR_c_301_n 0.00769046f $X=3.285 $Y=2.545 $X2=0
+ $Y2=0
cc_172 N_A_350_109#_M1003_g N_VPWR_c_295_n 0.0140911f $X=3.285 $Y=2.545 $X2=0
+ $Y2=0
cc_173 N_A_350_109#_c_233_n N_VPWR_c_295_n 0.021987f $X=2.13 $Y=2.19 $X2=0 $Y2=0
cc_174 N_A_350_109#_M1005_g X 0.0358729f $X=3.335 $Y=0.755 $X2=0 $Y2=0
cc_175 N_A_350_109#_c_234_n X 0.014089f $X=2.935 $Y=1.76 $X2=0 $Y2=0
cc_176 N_A_350_109#_c_229_n X 0.0390149f $X=3.1 $Y=1.34 $X2=0 $Y2=0
cc_177 N_A_350_109#_M1003_g X 0.015872f $X=3.285 $Y=2.545 $X2=0 $Y2=0
cc_178 N_A_350_109#_M1010_g N_X_c_330_n 5.77406e-19 $X=2.975 $Y=0.755 $X2=0
+ $Y2=0
cc_179 N_A_350_109#_M1005_g N_X_c_330_n 0.00825826f $X=3.335 $Y=0.755 $X2=0
+ $Y2=0
cc_180 N_A_350_109#_M1003_g X 0.00451956f $X=3.285 $Y=2.545 $X2=0 $Y2=0
cc_181 N_A_350_109#_c_231_n N_KAGND_c_349_n 0.00941356f $X=1.89 $Y=0.8 $X2=0
+ $Y2=0
cc_182 N_A_350_109#_c_231_n N_KAGND_c_350_n 0.0205125f $X=1.89 $Y=0.8 $X2=0
+ $Y2=0
cc_183 N_A_350_109#_M1010_g N_KAGND_c_351_n 0.0174483f $X=2.975 $Y=0.755 $X2=0
+ $Y2=0
cc_184 N_A_350_109#_M1005_g N_KAGND_c_351_n 0.00358937f $X=3.335 $Y=0.755 $X2=0
+ $Y2=0
cc_185 N_A_350_109#_c_229_n N_KAGND_c_351_n 0.0103695f $X=3.1 $Y=1.34 $X2=0
+ $Y2=0
cc_186 N_A_350_109#_c_231_n N_KAGND_c_351_n 0.00174654f $X=1.89 $Y=0.8 $X2=0
+ $Y2=0
cc_187 N_A_350_109#_M1004_d N_KAGND_c_352_n 6.62301e-19 $X=1.75 $Y=0.545 $X2=0
+ $Y2=0
cc_188 N_A_350_109#_M1005_g N_KAGND_c_352_n 0.00815779f $X=3.335 $Y=0.755 $X2=0
+ $Y2=0
cc_189 N_A_350_109#_c_228_n N_KAGND_c_352_n 5.27493e-19 $X=1.78 $Y=1.675 $X2=0
+ $Y2=0
cc_190 N_A_350_109#_c_229_n N_KAGND_c_352_n 0.00731488f $X=3.1 $Y=1.34 $X2=0
+ $Y2=0
cc_191 N_A_350_109#_c_231_n N_KAGND_c_352_n 0.0178133f $X=1.89 $Y=0.8 $X2=0
+ $Y2=0
cc_192 N_A_350_109#_M1005_g N_VGND_c_400_n 0.00293597f $X=3.335 $Y=0.755 $X2=0
+ $Y2=0
cc_193 N_A_350_109#_M1010_g N_VGND_c_401_n 6.46133e-19 $X=2.975 $Y=0.755 $X2=0
+ $Y2=0
cc_194 N_A_350_109#_M1005_g N_VGND_c_401_n 0.00441768f $X=3.335 $Y=0.755 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_301_n X 0.0220321f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_295_n X 0.0125808f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_297_n X 0.0684934f $X=3.02 $Y=2.19 $X2=0 $Y2=0
cc_198 N_X_c_330_n N_KAGND_c_351_n 0.0118897f $X=3.55 $Y=0.755 $X2=0 $Y2=0
cc_199 N_X_c_330_n N_KAGND_c_352_n 0.0320976f $X=3.55 $Y=0.755 $X2=0 $Y2=0
cc_200 N_X_c_330_n N_VGND_c_400_n 0.00142143f $X=3.55 $Y=0.755 $X2=0 $Y2=0
cc_201 N_X_c_330_n N_VGND_c_401_n 0.00876029f $X=3.55 $Y=0.755 $X2=0 $Y2=0
cc_202 A_114_109# N_KAGND_c_352_n 0.00225673f $X=0.57 $Y=0.545 $X2=2.94
+ $Y2=0.555
cc_203 N_KAGND_c_352_n A_272_109# 0.0051671f $X=2.94 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_204 N_KAGND_c_352_n A_452_109# 0.00225673f $X=2.94 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_205 N_KAGND_c_352_n A_610_109# 0.00227979f $X=2.94 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_206 N_KAGND_c_349_n N_VGND_c_400_n 0.0241654f $X=1.385 $Y=0.625 $X2=0 $Y2=0
cc_207 N_KAGND_c_352_n N_VGND_c_400_n 0.339561f $X=2.94 $Y=0.555 $X2=0 $Y2=0
cc_208 N_KAGND_c_349_n N_VGND_c_401_n 0.149645f $X=1.385 $Y=0.625 $X2=0 $Y2=0
cc_209 N_KAGND_c_352_n N_VGND_c_401_n 0.00737154f $X=2.94 $Y=0.555 $X2=0 $Y2=0
