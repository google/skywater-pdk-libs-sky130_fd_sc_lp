* File: sky130_fd_sc_lp__o22a_1.pex.spice
* Created: Wed Sep  2 10:19:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22A_1%A_80_21# 1 2 7 9 12 14 15 16 19 20 22 23 26
+ 28 30 32 38
r69 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.715
+ $Y=1.35 $X2=0.715 $Y2=1.35
r70 32 35 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.715 $Y=1.16
+ $X2=0.715 $Y2=1.35
r71 28 40 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.27 $Y=2.1 $X2=2.27
+ $Y2=2.015
r72 28 30 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=2.27 $Y=2.1
+ $X2=2.27 $Y2=2.775
r73 24 26 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=1.9 $Y=1.075
+ $X2=1.9 $Y2=0.93
r74 22 40 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.165 $Y=2.015
+ $X2=2.27 $Y2=2.015
r75 22 23 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.165 $Y=2.015 $X2=1.23
+ $Y2=2.015
r76 21 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=1.16
+ $X2=1.145 $Y2=1.16
r77 20 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.795 $Y=1.16
+ $X2=1.9 $Y2=1.075
r78 20 21 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.795 $Y=1.16
+ $X2=1.23 $Y2=1.16
r79 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=1.93
+ $X2=1.23 $Y2=2.015
r80 18 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.245
+ $X2=1.145 $Y2=1.16
r81 18 19 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.145 $Y=1.245
+ $X2=1.145 $Y2=1.93
r82 17 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=1.16
+ $X2=0.715 $Y2=1.16
r83 16 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=1.16
+ $X2=1.145 $Y2=1.16
r84 16 17 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.06 $Y=1.16
+ $X2=0.88 $Y2=1.16
r85 15 36 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.915 $Y=1.35
+ $X2=0.715 $Y2=1.35
r86 14 36 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.35
+ $X2=0.715 $Y2=1.35
r87 10 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.99 $Y=1.515
+ $X2=0.915 $Y2=1.35
r88 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.99 $Y=1.515
+ $X2=0.99 $Y2=2.465
r89 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.55 $Y2=1.35
r90 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
r91 2 40 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.835 $X2=2.27 $Y2=2.095
r92 2 30 400 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.835 $X2=2.27 $Y2=2.775
r93 1 26 182 $w=1.7e-07 $l=7.7086e-07 $layer=licon1_NDIFF $count=1 $X=1.74
+ $Y=0.235 $X2=1.9 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%B1 3 7 9 12 13
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.51
+ $X2=1.575 $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.51
+ $X2=1.575 $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=1.51 $X2=1.575 $Y2=1.51
r37 9 13 5.03179 $w=3.53e-07 $l=1.55e-07 $layer=LI1_cond $X=1.587 $Y=1.665
+ $X2=1.587 $Y2=1.51
r38 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.665 $Y=2.465
+ $X2=1.665 $Y2=1.675
r39 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.665 $Y=0.655
+ $X2=1.665 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%B2 3 7 9 12 13
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.51
+ $X2=2.145 $Y2=1.675
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.51
+ $X2=2.145 $Y2=1.345
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.145
+ $Y=1.51 $X2=2.145 $Y2=1.51
r39 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.145 $Y=1.665
+ $X2=2.145 $Y2=1.51
r40 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.115 $Y=0.655
+ $X2=2.115 $Y2=1.345
r41 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.055 $Y=2.465
+ $X2=2.055 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%A2 3 7 9 10 11 12 26 27
r37 26 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.51
+ $X2=2.74 $Y2=1.675
r38 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.51
+ $X2=2.74 $Y2=1.345
r39 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.51 $X2=2.74 $Y2=1.51
r40 11 12 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=2.405
+ $X2=2.88 $Y2=2.775
r41 10 11 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=2.035
+ $X2=2.88 $Y2=2.405
r42 9 10 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=2.035
r43 9 27 2.85219 $w=6.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=1.51
r44 7 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.65 $Y=2.465
+ $X2=2.65 $Y2=1.675
r45 3 28 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.65 $Y=0.655
+ $X2=2.65 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%A1 3 7 9 14 15
r24 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.46 $X2=3.55 $Y2=1.46
r25 11 14 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.22 $Y=1.46
+ $X2=3.55 $Y2=1.46
r26 9 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=1.46
r27 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.625
+ $X2=3.22 $Y2=1.46
r28 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.22 $Y=1.625 $X2=3.22
+ $Y2=2.465
r29 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.295
+ $X2=3.22 $Y2=1.46
r30 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.22 $Y=1.295 $X2=3.22
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%X 1 2 7 9 11 15 16 17 18 19 20 21 43
r24 41 43 2.64069 $w=2.08e-07 $l=5e-08 $layer=LI1_cond $X=0.26 $Y=1.985 $X2=0.26
+ $Y2=2.035
r25 20 21 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r26 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.9 $X2=0.26
+ $Y2=1.815
r27 19 41 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.9 $X2=0.26
+ $Y2=1.985
r28 19 20 18.6433 $w=2.08e-07 $l=3.53e-07 $layer=LI1_cond $X=0.26 $Y=2.052
+ $X2=0.26 $Y2=2.405
r29 19 43 0.897835 $w=2.08e-07 $l=1.7e-08 $layer=LI1_cond $X=0.26 $Y=2.052
+ $X2=0.26 $Y2=2.035
r30 18 30 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.815
r31 17 18 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r32 16 17 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.925
+ $X2=0.26 $Y2=1.295
r33 15 16 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.555
+ $X2=0.26 $Y2=0.925
r34 9 14 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=1.985
+ $X2=0.775 $Y2=1.9
r35 9 11 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.775 $Y=1.985
+ $X2=0.775 $Y2=2.66
r36 8 19 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.365 $Y=1.9 $X2=0.26
+ $Y2=1.9
r37 7 14 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.67 $Y=1.9 $X2=0.775
+ $Y2=1.9
r38 7 8 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.67 $Y=1.9 $X2=0.365
+ $Y2=1.9
r39 2 14 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.835 $X2=0.775 $Y2=1.98
r40 2 11 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.835 $X2=0.775 $Y2=2.66
r41 1 15 91 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%VPWR 1 2 9 11 13 17 19 24 33 37
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 25 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.205 $Y2=3.33
r49 25 27 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.31 $Y=3.33 $X2=1.68
+ $Y2=3.33
r50 24 36 3.61693 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.612 $Y2=3.33
r51 24 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 19 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=1.205 $Y2=3.33
r55 19 21 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r56 17 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 13 16 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=3.49 $Y=2.27
+ $X2=3.49 $Y2=2.95
r59 11 36 3.29826 $w=2.1e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.49 $Y=3.245
+ $X2=3.612 $Y2=3.33
r60 11 16 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.49 $Y=3.245
+ $X2=3.49 $Y2=2.95
r61 7 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=3.33
r62 7 9 33.5368 $w=2.08e-07 $l=6.35e-07 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=2.61
r63 2 16 400 $w=1.7e-07 $l=1.20857e-06 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.835 $X2=3.49 $Y2=2.95
r64 2 13 400 $w=1.7e-07 $l=5.23498e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.835 $X2=3.49 $Y2=2.27
r65 1 9 300 $w=1.7e-07 $l=8.42096e-07 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=1.835 $X2=1.205 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%VGND 1 2 9 13 16 17 18 20 30 31 34
r45 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r48 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 25 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.69
+ $Y2=0
r50 25 27 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=2.64 $Y2=0
r51 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r52 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 20 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.69
+ $Y2=0
r54 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r55 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r56 18 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.72
+ $Y2=0
r57 16 27 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.64
+ $Y2=0
r58 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.865
+ $Y2=0
r59 15 30 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.6
+ $Y2=0
r60 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.865
+ $Y2=0
r61 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0
r62 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0.38
r63 7 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r64 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r65 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=0.235 $X2=2.865 $Y2=0.38
r66 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_1%A_265_47# 1 2 3 12 14 15 16 17 20 23
r39 18 20 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=3.435 $Y=1.005
+ $X2=3.435 $Y2=0.59
r40 16 18 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.33 $Y=1.09
+ $X2=3.435 $Y2=1.005
r41 16 17 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.33 $Y=1.09
+ $X2=2.435 $Y2=1.09
r42 15 17 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.33 $Y=1.005
+ $X2=2.435 $Y2=1.09
r43 14 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.33 $Y=0.515
+ $X2=2.33 $Y2=0.43
r44 14 15 25.8788 $w=2.08e-07 $l=4.9e-07 $layer=LI1_cond $X=2.33 $Y=0.515
+ $X2=2.33 $Y2=1.005
r45 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0.43
+ $X2=1.45 $Y2=0.43
r46 12 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.225 $Y=0.43
+ $X2=2.33 $Y2=0.43
r47 12 13 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.225 $Y=0.43
+ $X2=1.615 $Y2=0.43
r48 3 20 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=3.295
+ $Y=0.235 $X2=3.435 $Y2=0.59
r49 2 25 91 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=2 $X=2.19
+ $Y=0.235 $X2=2.33 $Y2=0.51
r50 1 23 91 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=2 $X=1.325
+ $Y=0.235 $X2=1.45 $Y2=0.45
.ends

