* File: sky130_fd_sc_lp__nor4b_m.pxi.spice
* Created: Fri Aug 28 10:58:46 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4B_M%D_N N_D_N_M1008_g N_D_N_M1001_g N_D_N_c_78_n
+ N_D_N_c_83_n D_N D_N D_N D_N D_N N_D_N_c_80_n PM_SKY130_FD_SC_LP__NOR4B_M%D_N
x_PM_SKY130_FD_SC_LP__NOR4B_M%A N_A_c_123_n N_A_M1000_g N_A_c_128_n N_A_M1005_g
+ N_A_c_125_n N_A_c_131_n A A A A N_A_c_127_n PM_SKY130_FD_SC_LP__NOR4B_M%A
x_PM_SKY130_FD_SC_LP__NOR4B_M%B N_B_M1004_g N_B_M1006_g N_B_c_179_n N_B_c_184_n
+ B B B N_B_c_181_n PM_SKY130_FD_SC_LP__NOR4B_M%B
x_PM_SKY130_FD_SC_LP__NOR4B_M%C N_C_M1007_g N_C_M1009_g N_C_c_223_n N_C_c_228_n
+ C C C N_C_c_225_n PM_SKY130_FD_SC_LP__NOR4B_M%C
x_PM_SKY130_FD_SC_LP__NOR4B_M%A_33_68# N_A_33_68#_M1008_s N_A_33_68#_M1001_s
+ N_A_33_68#_M1003_g N_A_33_68#_c_267_n N_A_33_68#_M1002_g N_A_33_68#_c_274_n
+ N_A_33_68#_c_268_n N_A_33_68#_c_269_n N_A_33_68#_c_270_n N_A_33_68#_c_276_n
+ N_A_33_68#_c_277_n N_A_33_68#_c_278_n N_A_33_68#_c_279_n N_A_33_68#_c_271_n
+ N_A_33_68#_c_272_n N_A_33_68#_c_282_n PM_SKY130_FD_SC_LP__NOR4B_M%A_33_68#
x_PM_SKY130_FD_SC_LP__NOR4B_M%VPWR N_VPWR_M1001_d N_VPWR_c_343_n VPWR
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_342_n N_VPWR_c_347_n
+ PM_SKY130_FD_SC_LP__NOR4B_M%VPWR
x_PM_SKY130_FD_SC_LP__NOR4B_M%Y N_Y_M1000_d N_Y_M1009_d N_Y_M1003_d N_Y_c_368_n
+ N_Y_c_377_n N_Y_c_369_n N_Y_c_370_n N_Y_c_375_n N_Y_c_371_n Y Y Y Y
+ N_Y_c_374_n PM_SKY130_FD_SC_LP__NOR4B_M%Y
x_PM_SKY130_FD_SC_LP__NOR4B_M%VGND N_VGND_M1008_d N_VGND_M1004_d N_VGND_M1002_d
+ N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n N_VGND_c_422_n N_VGND_c_423_n
+ N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n
+ VGND N_VGND_c_429_n PM_SKY130_FD_SC_LP__NOR4B_M%VGND
cc_1 VNB N_D_N_M1008_g 0.0564138f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.55
cc_2 VNB N_D_N_c_78_n 5.7437e-19 $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.97
cc_3 VNB D_N 0.00667429f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_4 VNB N_D_N_c_80_n 0.0237104f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.615
cc_5 VNB N_A_c_123_n 0.0244923f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.55
cc_6 VNB N_A_M1000_g 0.0308844f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.647
cc_7 VNB N_A_c_125_n 0.00677758f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_8 VNB A 0.00365671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_127_n 0.0196867f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.555
cc_10 VNB N_B_M1004_g 0.0352761f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.55
cc_11 VNB N_B_c_179_n 0.0190398f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.97
cc_12 VNB B 9.23459e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_13 VNB N_B_c_181_n 0.0163122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C_M1009_g 0.0386934f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.12
cc_15 VNB N_C_c_223_n 0.0144619f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.97
cc_16 VNB C 0.00507986f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_17 VNB N_C_c_225_n 0.0154652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_33_68#_c_267_n 0.0212312f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.97
cc_19 VNB N_A_33_68#_c_268_n 0.0165164f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.615
cc_20 VNB N_A_33_68#_c_269_n 0.0369736f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.45
cc_21 VNB N_A_33_68#_c_270_n 0.0437087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_33_68#_c_271_n 0.0031683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_33_68#_c_272_n 0.00591511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_342_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_368_n 0.00138699f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.12
cc_26 VNB N_Y_c_369_n 0.0124347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_370_n 0.00445149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_371_n 0.032677f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.555
cc_29 VNB Y 0.0051332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 0.0114631f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.295
cc_31 VNB N_Y_c_374_n 0.0117734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_419_n 0.00783894f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.12
cc_33 VNB N_VGND_c_420_n 0.0071372f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_VGND_c_421_n 0.017987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_422_n 0.0307194f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.615
cc_36 VNB N_VGND_c_423_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.615
cc_37 VNB N_VGND_c_424_n 0.0197731f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.45
cc_38 VNB N_VGND_c_425_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.555
cc_39 VNB N_VGND_c_426_n 0.011849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_427_n 0.0190584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_428_n 0.0059043f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.925
cc_42 VNB N_VGND_c_429_n 0.214148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_D_N_M1001_g 0.0363376f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.69
cc_44 VPB N_D_N_c_78_n 0.0274778f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.97
cc_45 VPB N_D_N_c_83_n 0.0377756f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.12
cc_46 VPB D_N 0.00217992f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_47 VPB N_A_c_128_n 0.0197658f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.69
cc_48 VPB N_A_M1005_g 0.0206876f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.97
cc_49 VPB N_A_c_125_n 0.011289f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_50 VPB N_A_c_131_n 0.0243422f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_51 VPB A 0.00404516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_B_M1006_g 0.0375897f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.12
cc_53 VPB N_B_c_179_n 0.00402634f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.97
cc_54 VPB N_B_c_184_n 0.0164125f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.12
cc_55 VPB B 0.0034834f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_56 VPB N_C_M1007_g 0.034297f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.55
cc_57 VPB N_C_c_223_n 0.00672938f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.97
cc_58 VPB N_C_c_228_n 0.0154343f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.12
cc_59 VPB C 0.00582324f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_60 VPB N_A_33_68#_M1003_g 0.0231166f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.69
cc_61 VPB N_A_33_68#_c_274_n 0.0572151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_33_68#_c_270_n 0.0327048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_33_68#_c_276_n 0.00828804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_33_68#_c_277_n 0.0125645f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.295
cc_65 VPB N_A_33_68#_c_278_n 4.12885e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_33_68#_c_279_n 0.0421484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_33_68#_c_271_n 0.00347762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_33_68#_c_272_n 0.0109709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_33_68#_c_282_n 0.00184766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_343_n 0.0115409f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.97
cc_71 VPB N_VPWR_c_344_n 0.0333247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_345_n 0.0641679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_342_n 0.0897603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_347_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.615
cc_75 VPB N_Y_c_375_n 0.0162194f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.45
cc_76 VPB N_Y_c_371_n 0.0401446f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.555
cc_77 D_N N_A_c_123_n 0.00100798f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_78 N_D_N_c_80_n N_A_c_123_n 0.00880586f $X=0.66 $Y=1.615 $X2=0 $Y2=0
cc_79 N_D_N_M1008_g N_A_M1000_g 0.00788953f $X=0.505 $Y=0.55 $X2=0 $Y2=0
cc_80 D_N N_A_M1000_g 0.00433139f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_81 N_D_N_c_78_n N_A_c_128_n 0.00635652f $X=0.725 $Y=1.97 $X2=0 $Y2=0
cc_82 N_D_N_c_83_n N_A_c_128_n 0.0100552f $X=0.725 $Y=2.12 $X2=0 $Y2=0
cc_83 D_N N_A_c_128_n 3.75444e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_84 N_D_N_M1001_g N_A_M1005_g 0.0161732f $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_85 N_D_N_c_78_n N_A_c_125_n 0.00880586f $X=0.725 $Y=1.97 $X2=0 $Y2=0
cc_86 N_D_N_M1001_g N_A_c_131_n 0.0100552f $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_87 N_D_N_M1008_g A 9.20018e-19 $X=0.505 $Y=0.55 $X2=0 $Y2=0
cc_88 N_D_N_c_78_n A 0.00182063f $X=0.725 $Y=1.97 $X2=0 $Y2=0
cc_89 N_D_N_c_83_n A 0.00126998f $X=0.725 $Y=2.12 $X2=0 $Y2=0
cc_90 D_N A 0.0596368f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_91 N_D_N_c_80_n A 9.05006e-19 $X=0.66 $Y=1.615 $X2=0 $Y2=0
cc_92 N_D_N_M1008_g N_A_c_127_n 0.00838494f $X=0.505 $Y=0.55 $X2=0 $Y2=0
cc_93 D_N N_A_c_127_n 0.00354369f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_94 N_D_N_M1008_g N_A_33_68#_c_270_n 0.0345157f $X=0.505 $Y=0.55 $X2=0 $Y2=0
cc_95 N_D_N_M1001_g N_A_33_68#_c_270_n 0.00455994f $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_96 D_N N_A_33_68#_c_270_n 0.106561f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_97 N_D_N_c_83_n N_A_33_68#_c_276_n 0.00632964f $X=0.725 $Y=2.12 $X2=0 $Y2=0
cc_98 D_N N_A_33_68#_c_276_n 0.00371295f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_99 N_D_N_M1001_g N_A_33_68#_c_278_n 3.64605e-19 $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_100 N_D_N_M1001_g N_A_33_68#_c_279_n 0.0183435f $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_101 N_D_N_c_83_n N_A_33_68#_c_279_n 0.00116826f $X=0.725 $Y=2.12 $X2=0 $Y2=0
cc_102 N_D_N_c_83_n N_A_33_68#_c_282_n 0.00268778f $X=0.725 $Y=2.12 $X2=0 $Y2=0
cc_103 D_N N_A_33_68#_c_282_n 0.0148952f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_104 N_D_N_M1001_g N_VPWR_c_343_n 0.0130458f $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_105 N_D_N_M1001_g N_VPWR_c_344_n 0.00515352f $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_106 N_D_N_M1001_g N_VPWR_c_342_n 0.0051274f $X=0.945 $Y=2.69 $X2=0 $Y2=0
cc_107 D_N N_Y_c_377_n 2.71997e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_108 D_N N_VGND_M1008_d 0.00650377f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_109 N_D_N_M1008_g N_VGND_c_419_n 0.00480989f $X=0.505 $Y=0.55 $X2=0 $Y2=0
cc_110 D_N N_VGND_c_419_n 0.0129257f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_111 N_D_N_M1008_g N_VGND_c_422_n 0.00482212f $X=0.505 $Y=0.55 $X2=0 $Y2=0
cc_112 D_N N_VGND_c_422_n 0.00582308f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_113 N_D_N_M1008_g N_VGND_c_429_n 0.00989214f $X=0.505 $Y=0.55 $X2=0 $Y2=0
cc_114 D_N N_VGND_c_429_n 0.00776872f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A_M1000_g N_B_M1004_g 0.0266047f $X=1.305 $Y=0.55 $X2=0 $Y2=0
cc_116 A N_B_M1004_g 0.00119065f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_117 N_A_c_128_n N_B_M1006_g 0.00615206f $X=1.305 $Y=2.12 $X2=0 $Y2=0
cc_118 N_A_c_131_n N_B_M1006_g 0.0589111f $X=1.485 $Y=2.195 $X2=0 $Y2=0
cc_119 A N_B_M1006_g 2.16551e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_120 N_A_c_123_n N_B_c_179_n 0.0136749f $X=1.207 $Y=1.558 $X2=0 $Y2=0
cc_121 N_A_c_125_n N_B_c_184_n 0.0136749f $X=1.207 $Y=1.73 $X2=0 $Y2=0
cc_122 N_A_c_128_n B 0.0018829f $X=1.305 $Y=2.12 $X2=0 $Y2=0
cc_123 A B 0.0400828f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_124 N_A_c_127_n B 0.00242226f $X=1.2 $Y=1.225 $X2=0 $Y2=0
cc_125 A N_B_c_181_n 0.00203151f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_126 N_A_c_127_n N_B_c_181_n 0.0136749f $X=1.2 $Y=1.225 $X2=0 $Y2=0
cc_127 N_A_M1005_g N_A_33_68#_c_279_n 0.015719f $X=1.485 $Y=2.69 $X2=0 $Y2=0
cc_128 N_A_c_125_n N_A_33_68#_c_279_n 0.00254923f $X=1.207 $Y=1.73 $X2=0 $Y2=0
cc_129 N_A_c_131_n N_A_33_68#_c_279_n 0.00752682f $X=1.485 $Y=2.195 $X2=0 $Y2=0
cc_130 A N_A_33_68#_c_279_n 0.0133771f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_131 N_A_M1005_g N_VPWR_c_343_n 0.0106903f $X=1.485 $Y=2.69 $X2=0 $Y2=0
cc_132 N_A_M1005_g N_VPWR_c_345_n 0.00534427f $X=1.485 $Y=2.69 $X2=0 $Y2=0
cc_133 N_A_M1005_g N_VPWR_c_342_n 0.00526787f $X=1.485 $Y=2.69 $X2=0 $Y2=0
cc_134 N_A_M1000_g N_Y_c_377_n 0.00380822f $X=1.305 $Y=0.55 $X2=0 $Y2=0
cc_135 N_A_M1000_g Y 0.00488851f $X=1.305 $Y=0.55 $X2=0 $Y2=0
cc_136 A Y 0.0109476f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_137 N_A_M1000_g N_VGND_c_419_n 0.00353795f $X=1.305 $Y=0.55 $X2=0 $Y2=0
cc_138 A N_VGND_c_419_n 0.00470757f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_139 N_A_c_127_n N_VGND_c_419_n 0.00329125f $X=1.2 $Y=1.225 $X2=0 $Y2=0
cc_140 N_A_M1000_g N_VGND_c_424_n 0.00459209f $X=1.305 $Y=0.55 $X2=0 $Y2=0
cc_141 N_A_M1000_g N_VGND_c_429_n 0.00726139f $X=1.305 $Y=0.55 $X2=0 $Y2=0
cc_142 A N_VGND_c_429_n 0.00414425f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_143 N_B_M1006_g N_C_M1007_g 0.0279952f $X=1.845 $Y=2.69 $X2=0 $Y2=0
cc_144 N_B_M1004_g N_C_M1009_g 0.0263172f $X=1.735 $Y=0.55 $X2=0 $Y2=0
cc_145 N_B_c_181_n N_C_M1009_g 0.00245588f $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_146 N_B_c_179_n N_C_c_223_n 0.0279952f $X=1.755 $Y=1.715 $X2=0 $Y2=0
cc_147 N_B_c_184_n N_C_c_228_n 0.0279952f $X=1.755 $Y=1.88 $X2=0 $Y2=0
cc_148 B C 0.0549362f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_149 N_B_c_181_n C 0.00594205f $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_150 B N_C_c_225_n 8.7184e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_151 N_B_c_181_n N_C_c_225_n 0.0279952f $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_152 N_B_M1006_g N_A_33_68#_c_279_n 0.0134355f $X=1.845 $Y=2.69 $X2=0 $Y2=0
cc_153 N_B_c_184_n N_A_33_68#_c_279_n 8.90213e-19 $X=1.755 $Y=1.88 $X2=0 $Y2=0
cc_154 B N_A_33_68#_c_279_n 0.0191312f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B_M1006_g N_VPWR_c_345_n 0.00534427f $X=1.845 $Y=2.69 $X2=0 $Y2=0
cc_156 N_B_M1006_g N_VPWR_c_342_n 0.00526787f $X=1.845 $Y=2.69 $X2=0 $Y2=0
cc_157 N_B_M1004_g N_Y_c_377_n 0.0027064f $X=1.735 $Y=0.55 $X2=0 $Y2=0
cc_158 N_B_M1004_g N_Y_c_369_n 0.00906914f $X=1.735 $Y=0.55 $X2=0 $Y2=0
cc_159 B N_Y_c_369_n 0.0103733f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_160 N_B_c_181_n N_Y_c_369_n 0.00344999f $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_161 N_B_M1004_g Y 0.00638733f $X=1.735 $Y=0.55 $X2=0 $Y2=0
cc_162 B Y 0.00656098f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_B_c_181_n Y 7.16467e-19 $X=1.755 $Y=1.375 $X2=0 $Y2=0
cc_164 N_B_M1004_g N_VGND_c_420_n 0.00319486f $X=1.735 $Y=0.55 $X2=0 $Y2=0
cc_165 N_B_M1004_g N_VGND_c_424_n 0.00459209f $X=1.735 $Y=0.55 $X2=0 $Y2=0
cc_166 N_B_M1004_g N_VGND_c_429_n 0.0050194f $X=1.735 $Y=0.55 $X2=0 $Y2=0
cc_167 N_C_M1009_g N_A_33_68#_c_267_n 0.020009f $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_168 N_C_M1007_g N_A_33_68#_c_274_n 0.0626887f $X=2.205 $Y=2.69 $X2=0 $Y2=0
cc_169 N_C_c_228_n N_A_33_68#_c_274_n 0.00864322f $X=2.295 $Y=1.93 $X2=0 $Y2=0
cc_170 C N_A_33_68#_c_274_n 5.57077e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_171 N_C_M1009_g N_A_33_68#_c_269_n 0.00866438f $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_172 C N_A_33_68#_c_269_n 0.00312427f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_C_c_225_n N_A_33_68#_c_269_n 0.0209075f $X=2.295 $Y=1.425 $X2=0 $Y2=0
cc_174 N_C_M1007_g N_A_33_68#_c_279_n 0.0109915f $X=2.205 $Y=2.69 $X2=0 $Y2=0
cc_175 N_C_c_228_n N_A_33_68#_c_279_n 0.00313197f $X=2.295 $Y=1.93 $X2=0 $Y2=0
cc_176 C N_A_33_68#_c_279_n 0.0233202f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_177 N_C_M1007_g N_A_33_68#_c_271_n 0.00241403f $X=2.205 $Y=2.69 $X2=0 $Y2=0
cc_178 N_C_c_223_n N_A_33_68#_c_271_n 0.00187599f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_179 C N_A_33_68#_c_271_n 0.0364218f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_180 N_C_c_223_n N_A_33_68#_c_272_n 0.00864322f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_181 C N_A_33_68#_c_272_n 2.4997e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_C_M1007_g N_VPWR_c_345_n 0.00534427f $X=2.205 $Y=2.69 $X2=0 $Y2=0
cc_183 N_C_M1007_g N_VPWR_c_342_n 0.00526787f $X=2.205 $Y=2.69 $X2=0 $Y2=0
cc_184 N_C_M1009_g N_Y_c_368_n 0.00108434f $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_185 N_C_M1009_g N_Y_c_369_n 0.0124301f $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_186 C N_Y_c_369_n 0.0197047f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_187 N_C_c_225_n N_Y_c_369_n 4.43092e-19 $X=2.295 $Y=1.425 $X2=0 $Y2=0
cc_188 C N_Y_c_370_n 0.00197562f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_189 N_C_c_225_n N_Y_c_370_n 0.0036265f $X=2.295 $Y=1.425 $X2=0 $Y2=0
cc_190 N_C_M1009_g Y 5.66923e-19 $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_191 N_C_M1009_g N_VGND_c_420_n 0.00489553f $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_192 N_C_M1009_g N_VGND_c_421_n 7.35388e-19 $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_193 N_C_M1009_g N_VGND_c_427_n 0.00486513f $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_194 N_C_M1009_g N_VGND_c_429_n 0.00524419f $X=2.245 $Y=0.55 $X2=0 $Y2=0
cc_195 N_A_33_68#_c_279_n N_VPWR_c_343_n 0.0228571f $X=2.56 $Y=2.385 $X2=0 $Y2=0
cc_196 N_A_33_68#_c_278_n N_VPWR_c_344_n 0.00465601f $X=0.73 $Y=2.625 $X2=0
+ $Y2=0
cc_197 N_A_33_68#_M1003_g N_VPWR_c_345_n 0.00534427f $X=2.565 $Y=2.69 $X2=0
+ $Y2=0
cc_198 N_A_33_68#_M1003_g N_VPWR_c_342_n 0.00526787f $X=2.565 $Y=2.69 $X2=0
+ $Y2=0
cc_199 N_A_33_68#_c_276_n N_VPWR_c_342_n 0.00778021f $X=0.625 $Y=2.385 $X2=0
+ $Y2=0
cc_200 N_A_33_68#_c_277_n N_VPWR_c_342_n 0.00809722f $X=0.395 $Y=2.385 $X2=0
+ $Y2=0
cc_201 N_A_33_68#_c_278_n N_VPWR_c_342_n 0.00666966f $X=0.73 $Y=2.625 $X2=0
+ $Y2=0
cc_202 N_A_33_68#_c_279_n N_VPWR_c_342_n 0.0524978f $X=2.56 $Y=2.385 $X2=0 $Y2=0
cc_203 N_A_33_68#_c_267_n N_Y_c_368_n 0.00190976f $X=2.675 $Y=0.87 $X2=0 $Y2=0
cc_204 N_A_33_68#_M1003_g N_Y_c_375_n 0.0110708f $X=2.565 $Y=2.69 $X2=0 $Y2=0
cc_205 N_A_33_68#_c_274_n N_Y_c_375_n 0.00355248f $X=2.835 $Y=2.17 $X2=0 $Y2=0
cc_206 N_A_33_68#_c_279_n N_Y_c_375_n 7.87385e-19 $X=2.56 $Y=2.385 $X2=0 $Y2=0
cc_207 N_A_33_68#_M1003_g N_Y_c_371_n 0.00151865f $X=2.565 $Y=2.69 $X2=0 $Y2=0
cc_208 N_A_33_68#_c_268_n N_Y_c_371_n 0.0200811f $X=2.775 $Y=0.945 $X2=0 $Y2=0
cc_209 N_A_33_68#_c_279_n N_Y_c_371_n 0.00891337f $X=2.56 $Y=2.385 $X2=0 $Y2=0
cc_210 N_A_33_68#_c_271_n N_Y_c_371_n 0.0469904f $X=2.835 $Y=1.815 $X2=0 $Y2=0
cc_211 N_A_33_68#_c_272_n N_Y_c_371_n 0.0167063f $X=2.835 $Y=1.815 $X2=0 $Y2=0
cc_212 N_A_33_68#_c_267_n N_Y_c_374_n 0.00468185f $X=2.675 $Y=0.87 $X2=0 $Y2=0
cc_213 N_A_33_68#_c_268_n N_Y_c_374_n 0.0152142f $X=2.775 $Y=0.945 $X2=0 $Y2=0
cc_214 N_A_33_68#_c_271_n N_Y_c_374_n 0.00990519f $X=2.835 $Y=1.815 $X2=0 $Y2=0
cc_215 N_A_33_68#_c_272_n N_Y_c_374_n 0.00241776f $X=2.835 $Y=1.815 $X2=0 $Y2=0
cc_216 N_A_33_68#_c_267_n N_VGND_c_421_n 0.00942097f $X=2.675 $Y=0.87 $X2=0
+ $Y2=0
cc_217 N_A_33_68#_c_268_n N_VGND_c_421_n 4.98678e-19 $X=2.775 $Y=0.945 $X2=0
+ $Y2=0
cc_218 N_A_33_68#_c_270_n N_VGND_c_422_n 0.00608118f $X=0.29 $Y=0.615 $X2=0
+ $Y2=0
cc_219 N_A_33_68#_c_267_n N_VGND_c_427_n 0.0040395f $X=2.675 $Y=0.87 $X2=0 $Y2=0
cc_220 N_A_33_68#_c_267_n N_VGND_c_429_n 0.00404872f $X=2.675 $Y=0.87 $X2=0
+ $Y2=0
cc_221 N_A_33_68#_c_270_n N_VGND_c_429_n 0.00720343f $X=0.29 $Y=0.615 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_345_n N_Y_c_375_n 0.00922534f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_342_n N_Y_c_375_n 0.0116827f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_224 N_Y_c_369_n N_VGND_c_420_n 0.0153318f $X=2.355 $Y=0.925 $X2=0 $Y2=0
cc_225 N_Y_c_374_n N_VGND_c_421_n 0.0172791f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_226 N_Y_c_377_n N_VGND_c_424_n 0.00789072f $X=1.6 $Y=0.555 $X2=0 $Y2=0
cc_227 N_Y_c_368_n N_VGND_c_427_n 0.00538635f $X=2.46 $Y=0.615 $X2=0 $Y2=0
cc_228 N_Y_c_368_n N_VGND_c_429_n 0.00645427f $X=2.46 $Y=0.615 $X2=0 $Y2=0
cc_229 N_Y_c_377_n N_VGND_c_429_n 0.0106694f $X=1.6 $Y=0.555 $X2=0 $Y2=0
cc_230 N_Y_c_369_n N_VGND_c_429_n 0.014666f $X=2.355 $Y=0.925 $X2=0 $Y2=0
cc_231 Y N_VGND_c_429_n 0.00670311f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_232 N_Y_c_374_n N_VGND_c_429_n 0.00815222f $X=3.1 $Y=0.925 $X2=0 $Y2=0
