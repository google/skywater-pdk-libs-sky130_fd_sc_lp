* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 VGND D a_437_144# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_547_167# a_437_144# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR D a_437_144# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_955_271# a_630_167# a_1211_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND a_955_271# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_207_40# a_112_70# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_955_271# a_625_377# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND GATE_N a_112_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_955_271# a_1394_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VGND a_955_271# a_716_167# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_207_40# a_112_70# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_630_167# a_207_40# a_813_377# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_813_377# a_437_144# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VPWR a_955_271# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_547_167# a_112_70# a_630_167# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Q_N a_1394_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VGND a_955_271# a_1394_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_955_271# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR GATE_N a_112_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VPWR a_630_167# a_955_271# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_1211_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_625_377# a_112_70# a_630_167# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 Q_N a_1394_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_630_167# a_207_40# a_716_167# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
