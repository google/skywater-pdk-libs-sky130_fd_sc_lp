* File: sky130_fd_sc_lp__dlrbn_2.pex.spice
* Created: Wed Sep  2 09:46:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRBN_2%GATE_N 2 5 8 10 11 12 13 14 20 22
c31 20 0 6.25322e-20 $X=0.385 $Y=1.415
r32 20 22 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.415
+ $X2=0.407 $Y2=1.25
r33 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.415 $X2=0.385 $Y2=1.415
r34 13 14 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=2.035
+ $X2=0.277 $Y2=2.405
r35 12 13 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=2.035
r36 12 21 7.4834 $w=3.83e-07 $l=2.5e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.415
r37 11 21 3.59203 $w=3.83e-07 $l=1.2e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.415
r38 8 10 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.52 $Y=2.685
+ $X2=0.52 $Y2=1.92
r39 5 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.49 $Y=0.93 $X2=0.49
+ $Y2=1.25
r40 2 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.407 $Y=1.733
+ $X2=0.407 $Y2=1.92
r41 1 20 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.437
+ $X2=0.407 $Y2=1.415
r42 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.407 $Y=1.437
+ $X2=0.407 $Y2=1.733
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_113_144# 1 2 7 9 12 14 18 20 24 26 27 28
+ 30 34 35 37 41 48 55
c103 41 0 1.15562e-19 $X=0.705 $Y=0.865
c104 7 0 2.29586e-20 $X=1.455 $Y=1.25
r105 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.415 $X2=0.97 $Y2=1.415
r106 46 48 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.77 $Y=1.415 $X2=0.97
+ $Y2=1.415
r107 44 46 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=0.73 $Y=1.415 $X2=0.77
+ $Y2=1.415
r108 41 43 8.97179 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=0.865
+ $X2=0.715 $Y2=1.03
r109 38 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=2.94
+ $X2=1.52 $Y2=2.94
r110 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.355
+ $Y=2.94 $X2=1.355 $Y2=2.94
r111 35 37 17.4787 $w=2.98e-07 $l=4.55e-07 $layer=LI1_cond $X=0.9 $Y=2.925
+ $X2=1.355 $Y2=2.925
r112 32 35 6.86182 $w=3e-07 $l=2.04939e-07 $layer=LI1_cond $X=0.77 $Y=2.775
+ $X2=0.9 $Y2=2.925
r113 32 34 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.77 $Y=2.775
+ $X2=0.77 $Y2=2.52
r114 31 46 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.58
+ $X2=0.77 $Y2=1.415
r115 31 34 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=0.77 $Y=1.58
+ $X2=0.77 $Y2=2.52
r116 30 44 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=1.25
+ $X2=0.73 $Y2=1.415
r117 30 43 13.5556 $w=1.78e-07 $l=2.2e-07 $layer=LI1_cond $X=0.73 $Y=1.25
+ $X2=0.73 $Y2=1.03
r118 26 49 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.38 $Y=1.415
+ $X2=0.97 $Y2=1.415
r119 26 27 5.03009 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.38 $Y=1.415
+ $X2=1.475 $Y2=1.415
r120 22 24 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.37 $Y=2.805
+ $X2=3.37 $Y2=2.005
r121 21 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=2.88
+ $X2=2.88 $Y2=2.88
r122 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.295 $Y=2.88
+ $X2=3.37 $Y2=2.805
r123 20 21 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.295 $Y=2.88
+ $X2=2.955 $Y2=2.88
r124 16 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.88 $Y=2.805
+ $X2=2.88 $Y2=2.88
r125 16 18 933.234 $w=1.5e-07 $l=1.82e-06 $layer=POLY_cond $X=2.88 $Y=2.805
+ $X2=2.88 $Y2=0.985
r126 14 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.805 $Y=2.88
+ $X2=2.88 $Y2=2.88
r127 14 55 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=2.805 $Y=2.88
+ $X2=1.52 $Y2=2.88
r128 10 27 37.0704 $w=1.5e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.495 $Y=1.58
+ $X2=1.475 $Y2=1.415
r129 10 12 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.495 $Y=1.58
+ $X2=1.495 $Y2=2.115
r130 7 27 37.0704 $w=1.5e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.455 $Y=1.25
+ $X2=1.475 $Y2=1.415
r131 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.455 $Y=1.25
+ $X2=1.455 $Y2=0.93
r132 2 34 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.365 $X2=0.735 $Y2=2.52
r133 1 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.72 $X2=0.705 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%D 1 3 6 8 9 17
c34 1 0 2.89292e-20 $X=1.885 $Y=1.25
r35 15 17 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.945 $Y=1.415
+ $X2=2.08 $Y2=1.415
r36 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.945
+ $Y=1.415 $X2=1.945 $Y2=1.415
r37 12 15 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.885 $Y=1.415
+ $X2=1.945 $Y2=1.415
r38 9 16 6.57186 $w=4.53e-07 $l=2.5e-07 $layer=LI1_cond $X=1.802 $Y=1.665
+ $X2=1.802 $Y2=1.415
r39 8 16 3.15449 $w=4.53e-07 $l=1.2e-07 $layer=LI1_cond $X=1.802 $Y=1.295
+ $X2=1.802 $Y2=1.415
r40 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.58
+ $X2=2.08 $Y2=1.415
r41 4 6 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.08 $Y=1.58 $X2=2.08
+ $Y2=2.115
r42 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.25
+ $X2=1.885 $Y2=1.415
r43 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.885 $Y=1.25
+ $X2=1.885 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_162_40# 1 2 7 12 13 14 17 19 20 21 23 34
+ 36 37
c81 37 0 1.15562e-19 $X=0.975 $Y=0.275
c82 36 0 9.14615e-20 $X=1.26 $Y=1.775
c83 19 0 2.29586e-20 $X=1.24 $Y=0.45
r84 35 36 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.32 $Y=1.08
+ $X2=1.32 $Y2=1.775
r85 34 35 7.93834 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.24 $Y=0.93
+ $X2=1.24 $Y2=1.08
r86 29 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.975 $Y=0.365
+ $X2=0.975 $Y2=0.275
r87 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=0.365 $X2=0.975 $Y2=0.365
r88 21 36 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.26 $Y=1.92
+ $X2=1.26 $Y2=1.775
r89 21 23 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=1.26 $Y=1.92 $X2=1.26
+ $Y2=1.94
r90 20 34 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.24 $Y=0.915
+ $X2=1.24 $Y2=0.93
r91 19 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.24 $Y=0.365
+ $X2=0.975 $Y2=0.365
r92 19 20 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.24 $Y=0.45
+ $X2=1.24 $Y2=0.915
r93 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.895 $Y=1.455
+ $X2=3.895 $Y2=2.115
r94 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.82 $Y=1.38
+ $X2=3.895 $Y2=1.455
r95 13 14 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.82 $Y=1.38
+ $X2=3.385 $Y2=1.38
r96 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.31 $Y=1.305
+ $X2=3.385 $Y2=1.38
r97 10 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.31 $Y=1.305
+ $X2=3.31 $Y2=0.985
r98 9 12 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.31 $Y=0.35
+ $X2=3.31 $Y2=0.985
r99 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=0.275
+ $X2=0.975 $Y2=0.275
r100 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.235 $Y=0.275
+ $X2=3.31 $Y2=0.35
r101 7 8 1074.24 $w=1.5e-07 $l=2.095e-06 $layer=POLY_cond $X=3.235 $Y=0.275
+ $X2=1.14 $Y2=0.275
r102 2 23 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.155
+ $Y=1.795 $X2=1.28 $Y2=1.94
r103 1 34 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.72 $X2=1.24 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_392_144# 1 2 8 9 10 13 15 17 19 21 23 26
+ 28 29 31 32 38
c90 10 0 1.75139e-19 $X=3.955 $Y=1.01
r91 37 38 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.29 $Y=0.87
+ $X2=2.295 $Y2=0.87
r92 35 37 6.44012 $w=3.38e-07 $l=1.9e-07 $layer=LI1_cond $X=2.1 $Y=0.87 $X2=2.29
+ $Y2=0.87
r93 32 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=0.35
+ $X2=3.79 $Y2=0.515
r94 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.79
+ $Y=0.35 $X2=3.79 $Y2=0.35
r95 29 31 82.3062 $w=1.88e-07 $l=1.41e-06 $layer=LI1_cond $X=2.38 $Y=0.35
+ $X2=3.79 $Y2=0.35
r96 28 38 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.295 $Y=0.7
+ $X2=2.295 $Y2=0.87
r97 27 29 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.295 $Y=0.445
+ $X2=2.38 $Y2=0.35
r98 27 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.295 $Y=0.445
+ $X2=2.295 $Y2=0.7
r99 26 41 8.65715 $w=2.97e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.29 $Y=1.775
+ $X2=2.295 $Y2=1.94
r100 25 37 4.46199 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=2.29 $Y=1.04
+ $X2=2.29 $Y2=0.87
r101 25 26 45.2879 $w=1.78e-07 $l=7.35e-07 $layer=LI1_cond $X=2.29 $Y=1.04
+ $X2=2.29 $Y2=1.775
r102 21 41 5.5092 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=2.295 $Y=2.085
+ $X2=2.295 $Y2=1.94
r103 21 23 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.295 $Y=2.085
+ $X2=2.295 $Y2=2.28
r104 18 19 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.255 $Y=1.01
+ $X2=4.425 $Y2=1.01
r105 15 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.425 $Y=0.935
+ $X2=4.425 $Y2=1.01
r106 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.425 $Y=0.935
+ $X2=4.425 $Y2=0.615
r107 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.255 $Y=1.085
+ $X2=4.255 $Y2=1.01
r108 11 13 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=4.255 $Y=1.085
+ $X2=4.255 $Y2=2.115
r109 9 18 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=1.01
+ $X2=4.255 $Y2=1.01
r110 9 10 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.18 $Y=1.01
+ $X2=3.955 $Y2=1.01
r111 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.88 $Y=0.935
+ $X2=3.955 $Y2=1.01
r112 8 44 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.88 $Y=0.935
+ $X2=3.88 $Y2=0.515
r113 2 41 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.795 $X2=2.295 $Y2=1.94
r114 2 23 600 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.795 $X2=2.295 $Y2=2.28
r115 1 35 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.72 $X2=2.1 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_942_252# 1 2 9 13 17 21 25 29 33 37 39 44
+ 45 46 49 53 56 57 58 61 63 64 67 68 70 72
c147 70 0 1.88466e-20 $X=5.6 $Y=1.465
c148 56 0 7.75143e-20 $X=5.65 $Y=2.325
c149 29 0 2.61412e-19 $X=7.175 $Y=2.465
r150 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.49 $X2=7.31 $Y2=1.49
r151 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.99
+ $Y=1.49 $X2=7.99 $Y2=1.49
r152 65 74 5.07179 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=7.58 $Y=1.49
+ $X2=7.362 $Y2=1.49
r153 65 67 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.58 $Y=1.49
+ $X2=7.99 $Y2=1.49
r154 63 74 2.90814 $w=3.55e-07 $l=1.03078e-07 $layer=LI1_cond $X=7.402 $Y=1.575
+ $X2=7.362 $Y2=1.49
r155 63 64 24.3474 $w=3.53e-07 $l=7.5e-07 $layer=LI1_cond $X=7.402 $Y=1.575
+ $X2=7.402 $Y2=2.325
r156 62 72 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.175 $Y=2.41
+ $X2=6.055 $Y2=2.41
r157 61 64 7.97992 $w=1.7e-07 $l=2.15346e-07 $layer=LI1_cond $X=7.225 $Y=2.41
+ $X2=7.402 $Y2=2.325
r158 61 62 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=7.225 $Y=2.41
+ $X2=6.175 $Y2=2.41
r159 57 72 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.935 $Y=2.41
+ $X2=6.055 $Y2=2.41
r160 57 58 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.935 $Y=2.41
+ $X2=5.735 $Y2=2.41
r161 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.65 $Y=2.325
+ $X2=5.735 $Y2=2.41
r162 55 70 6.28297 $w=2.2e-07 $l=1.63095e-07 $layer=LI1_cond $X=5.65 $Y=1.605
+ $X2=5.6 $Y2=1.465
r163 55 56 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.65 $Y=1.605
+ $X2=5.65 $Y2=2.325
r164 51 70 6.28297 $w=2.2e-07 $l=1.4e-07 $layer=LI1_cond $X=5.6 $Y=1.325 $X2=5.6
+ $Y2=1.465
r165 51 53 37.5611 $w=2.68e-07 $l=8.8e-07 $layer=LI1_cond $X=5.6 $Y=1.325
+ $X2=5.6 $Y2=0.445
r166 49 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.425
+ $X2=4.875 $Y2=1.59
r167 49 80 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.425
+ $X2=4.875 $Y2=1.26
r168 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.425 $X2=4.875 $Y2=1.425
r169 46 70 0.490351 $w=2.8e-07 $l=1.35e-07 $layer=LI1_cond $X=5.465 $Y=1.465
+ $X2=5.6 $Y2=1.465
r170 46 48 24.2836 $w=2.78e-07 $l=5.9e-07 $layer=LI1_cond $X=5.465 $Y=1.465
+ $X2=4.875 $Y2=1.465
r171 44 75 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=7.625 $Y=1.49
+ $X2=7.31 $Y2=1.49
r172 44 45 4.10278 $w=3.3e-07 $l=8.2e-08 $layer=POLY_cond $X=7.625 $Y=1.49
+ $X2=7.707 $Y2=1.49
r173 43 68 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.79 $Y=1.49 $X2=7.99
+ $Y2=1.49
r174 43 45 4.10278 $w=3.3e-07 $l=8.3e-08 $layer=POLY_cond $X=7.79 $Y=1.49
+ $X2=7.707 $Y2=1.49
r175 40 42 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.745 $Y=1.49
+ $X2=7.175 $Y2=1.49
r176 39 75 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=7.25 $Y=1.49 $X2=7.31
+ $Y2=1.49
r177 39 42 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.25 $Y=1.49
+ $X2=7.175 $Y2=1.49
r178 35 45 22.6206 $w=1.5e-07 $l=1.68953e-07 $layer=POLY_cond $X=7.715 $Y=1.325
+ $X2=7.707 $Y2=1.49
r179 35 37 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.715 $Y=1.325
+ $X2=7.715 $Y2=0.93
r180 31 45 22.6206 $w=1.5e-07 $l=1.68464e-07 $layer=POLY_cond $X=7.7 $Y=1.655
+ $X2=7.707 $Y2=1.49
r181 31 33 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.7 $Y=1.655 $X2=7.7
+ $Y2=2.155
r182 27 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.175 $Y=1.655
+ $X2=7.175 $Y2=1.49
r183 27 29 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.175 $Y=1.655
+ $X2=7.175 $Y2=2.465
r184 23 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.175 $Y=1.325
+ $X2=7.175 $Y2=1.49
r185 23 25 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=7.175 $Y=1.325
+ $X2=7.175 $Y2=0.72
r186 19 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.745 $Y=1.655
+ $X2=6.745 $Y2=1.49
r187 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.745 $Y=1.655
+ $X2=6.745 $Y2=2.465
r188 15 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.745 $Y=1.325
+ $X2=6.745 $Y2=1.49
r189 15 17 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=6.745 $Y=1.325
+ $X2=6.745 $Y2=0.72
r190 13 80 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.855 $Y=0.615
+ $X2=4.855 $Y2=1.26
r191 9 81 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.785 $Y=2.005
+ $X2=4.785 $Y2=1.59
r192 2 72 300 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=2 $X=5.92
+ $Y=1.835 $X2=6.06 $Y2=2.49
r193 1 53 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.505
+ $Y=0.3 $X2=5.63 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_591_155# 1 2 7 10 11 12 15 17 19 20 22 23
+ 24 25 27 31 32 39
c101 27 0 7.7762e-20 $X=3.095 $Y=1.07
r102 39 40 8.67082 $w=4.01e-07 $l=2.85e-07 $layer=LI1_cond $X=3.68 $Y=2.355
+ $X2=3.965 $Y2=2.355
r103 32 43 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.965 $Y=2.94
+ $X2=3.965 $Y2=3.03
r104 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.965
+ $Y=2.94 $X2=3.965 $Y2=2.94
r105 29 40 1.88052 $w=3.3e-07 $l=2.4e-07 $layer=LI1_cond $X=3.965 $Y=2.595
+ $X2=3.965 $Y2=2.355
r106 29 31 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.965 $Y=2.595
+ $X2=3.965 $Y2=2.94
r107 25 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.095 $Y=1.51
+ $X2=2.785 $Y2=1.51
r108 25 27 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.095 $Y=1.425
+ $X2=3.095 $Y2=1.07
r109 23 39 5.68006 $w=4.01e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.515 $Y=2.44
+ $X2=3.68 $Y2=2.355
r110 23 24 23.9782 $w=3.08e-07 $l=6.45e-07 $layer=LI1_cond $X=3.515 $Y=2.44
+ $X2=2.87 $Y2=2.44
r111 22 24 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.785 $Y=2.285
+ $X2=2.87 $Y2=2.44
r112 21 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.595
+ $X2=2.785 $Y2=1.51
r113 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.785 $Y=1.595
+ $X2=2.785 $Y2=2.285
r114 17 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.845 $Y=1.725
+ $X2=5.845 $Y2=1.65
r115 17 19 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.845 $Y=1.725
+ $X2=5.845 $Y2=2.465
r116 13 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.845 $Y=1.575
+ $X2=5.845 $Y2=1.65
r117 13 15 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=5.845 $Y=1.575
+ $X2=5.845 $Y2=0.72
r118 11 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.77 $Y=1.65
+ $X2=5.845 $Y2=1.65
r119 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.77 $Y=1.65
+ $X2=5.43 $Y2=1.65
r120 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.355 $Y=1.725
+ $X2=5.43 $Y2=1.65
r121 9 10 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=5.355 $Y=1.725
+ $X2=5.355 $Y2=2.955
r122 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=3.03
+ $X2=3.965 $Y2=3.03
r123 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.28 $Y=3.03
+ $X2=5.355 $Y2=2.955
r124 7 8 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=5.28 $Y=3.03
+ $X2=4.13 $Y2=3.03
r125 2 39 600 $w=1.7e-07 $l=5.29622e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.795 $X2=3.68 $Y2=2.22
r126 1 27 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.775 $X2=3.095 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%RESET_B 3 6 8 9 10 21 23
c37 23 0 2.67944e-20 $X=6.295 $Y=1.25
c38 21 0 3.25769e-21 $X=6.295 $Y=1.415
c39 6 0 9.31032e-20 $X=6.275 $Y=2.465
r40 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=1.415
+ $X2=6.295 $Y2=1.58
r41 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=1.415
+ $X2=6.295 $Y2=1.25
r42 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.295
+ $Y=1.415 $X2=6.295 $Y2=1.415
r43 9 10 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=6.27 $Y=1.665
+ $X2=6.27 $Y2=2.035
r44 9 22 4.21154 $w=7.08e-07 $l=2.5e-07 $layer=LI1_cond $X=6.27 $Y=1.665
+ $X2=6.27 $Y2=1.415
r45 8 22 2.02154 $w=7.08e-07 $l=1.2e-07 $layer=LI1_cond $X=6.27 $Y=1.295
+ $X2=6.27 $Y2=1.415
r46 6 24 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=6.275 $Y=2.465
+ $X2=6.275 $Y2=1.58
r47 3 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.205 $Y=0.72
+ $X2=6.205 $Y2=1.25
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_1555_367# 1 2 9 13 15 19 23 25 28 30 34 35
+ 39 41
c65 35 0 1.16002e-19 $X=8.02 $Y=1.84
r66 41 42 32.8921 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=8.562 $Y=1.385
+ $X2=8.562 $Y2=1.31
r67 40 44 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=8.562 $Y=1.475
+ $X2=8.562 $Y2=1.64
r68 40 41 12.6719 $w=3.95e-07 $l=9e-08 $layer=POLY_cond $X=8.562 $Y=1.475
+ $X2=8.562 $Y2=1.385
r69 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.53
+ $Y=1.475 $X2=8.53 $Y2=1.475
r70 37 39 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=8.49 $Y=1.755
+ $X2=8.49 $Y2=1.475
r71 36 39 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=8.49 $Y=1.115
+ $X2=8.49 $Y2=1.475
r72 34 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.365 $Y=1.84
+ $X2=8.49 $Y2=1.755
r73 34 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.365 $Y=1.84
+ $X2=8.02 $Y2=1.84
r74 30 36 6.8319 $w=2.3e-07 $l=1.73205e-07 $layer=LI1_cond $X=8.365 $Y=1
+ $X2=8.49 $Y2=1.115
r75 30 32 21.7962 $w=2.28e-07 $l=4.35e-07 $layer=LI1_cond $X=8.365 $Y=1 $X2=7.93
+ $Y2=1
r76 26 35 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.885 $Y=1.925
+ $X2=8.02 $Y2=1.84
r77 26 28 2.34757 $w=2.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.885 $Y=1.925
+ $X2=7.885 $Y2=1.98
r78 21 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.115 $Y=1.46
+ $X2=9.115 $Y2=1.385
r79 21 23 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=9.115 $Y=1.46
+ $X2=9.115 $Y2=2.465
r80 17 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.115 $Y=1.31
+ $X2=9.115 $Y2=1.385
r81 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=9.115 $Y=1.31
+ $X2=9.115 $Y2=0.69
r82 16 41 25.5547 $w=1.5e-07 $l=1.98e-07 $layer=POLY_cond $X=8.76 $Y=1.385
+ $X2=8.562 $Y2=1.385
r83 15 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.04 $Y=1.385
+ $X2=9.115 $Y2=1.385
r84 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.04 $Y=1.385
+ $X2=8.76 $Y2=1.385
r85 13 44 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=8.685 $Y=2.465
+ $X2=8.685 $Y2=1.64
r86 9 42 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.685 $Y=0.69
+ $X2=8.685 $Y2=1.31
r87 2 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.775
+ $Y=1.835 $X2=7.915 $Y2=1.98
r88 1 32 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=7.79
+ $Y=0.72 $X2=7.93 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 43 47 51
+ 55 57 62 63 65 66 67 76 87 91 96 101 110 113 116 119 123
r126 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r127 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r128 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r129 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r130 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 105 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r133 105 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r134 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r135 102 119 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.465 $Y2=3.33
r136 102 104 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.88 $Y2=3.33
r137 101 122 4.38699 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=9.205 $Y=3.33
+ $X2=9.402 $Y2=3.33
r138 101 104 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=3.33
+ $X2=8.88 $Y2=3.33
r139 100 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r140 100 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r141 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r142 97 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.555 $Y=3.33
+ $X2=7.39 $Y2=3.33
r143 97 99 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.555 $Y=3.33
+ $X2=7.92 $Y2=3.33
r144 96 119 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.305 $Y=3.33
+ $X2=8.465 $Y2=3.33
r145 96 99 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.305 $Y=3.33
+ $X2=7.92 $Y2=3.33
r146 95 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r147 95 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r148 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 92 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.51 $Y2=3.33
r150 92 94 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.96 $Y2=3.33
r151 91 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.225 $Y=3.33
+ $X2=7.39 $Y2=3.33
r152 91 94 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.225 $Y=3.33
+ $X2=6.96 $Y2=3.33
r153 90 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r154 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r155 87 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.345 $Y=3.33
+ $X2=6.51 $Y2=3.33
r156 87 89 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.345 $Y=3.33 $X2=6
+ $Y2=3.33
r157 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r158 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r159 83 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=3.33
+ $X2=4.475 $Y2=3.33
r160 83 85 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=4.64 $Y=3.33
+ $X2=5.52 $Y2=3.33
r161 82 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r162 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r163 79 82 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r164 78 81 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r165 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r166 76 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=3.33
+ $X2=4.475 $Y2=3.33
r167 76 81 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.31 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 75 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r169 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r170 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r171 72 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r172 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r173 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 69 107 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.235 $Y2=3.33
r175 69 71 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.72 $Y2=3.33
r176 67 86 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r177 67 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r178 65 85 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.525 $Y=3.33
+ $X2=5.52 $Y2=3.33
r179 65 66 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.525 $Y=3.33
+ $X2=5.645 $Y2=3.33
r180 64 89 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=6 $Y2=3.33
r181 64 66 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.645 $Y2=3.33
r182 62 74 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.69 $Y=3.33
+ $X2=1.68 $Y2=3.33
r183 62 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.69 $Y=3.33
+ $X2=1.815 $Y2=3.33
r184 61 78 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.16 $Y2=3.33
r185 61 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.815 $Y2=3.33
r186 57 60 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=9.35 $Y=1.98
+ $X2=9.35 $Y2=2.95
r187 55 122 3.05085 $w=2.9e-07 $l=1.07912e-07 $layer=LI1_cond $X=9.35 $Y=3.245
+ $X2=9.402 $Y2=3.33
r188 55 60 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=9.35 $Y=3.245
+ $X2=9.35 $Y2=2.95
r189 51 54 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=8.465 $Y=2.27
+ $X2=8.465 $Y2=2.95
r190 49 119 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=3.33
r191 49 54 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=2.95
r192 45 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=3.33
r193 45 47 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=2.77
r194 41 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.51 $Y=3.245
+ $X2=6.51 $Y2=3.33
r195 41 43 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=6.51 $Y=3.245
+ $X2=6.51 $Y2=2.77
r196 37 66 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=3.33
r197 37 39 19.9277 $w=2.38e-07 $l=4.15e-07 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=2.83
r198 33 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=3.245
+ $X2=4.475 $Y2=3.33
r199 33 35 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=4.475 $Y=3.245
+ $X2=4.475 $Y2=2.245
r200 29 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=3.245
+ $X2=1.815 $Y2=3.33
r201 29 31 53.4734 $w=2.48e-07 $l=1.16e-06 $layer=LI1_cond $X=1.815 $Y=3.245
+ $X2=1.815 $Y2=2.085
r202 25 107 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.235 $Y2=3.33
r203 25 27 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.305 $Y2=2.785
r204 8 60 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.835 $X2=9.33 $Y2=2.95
r205 8 57 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.835 $X2=9.33 $Y2=1.98
r206 7 54 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=8.345
+ $Y=1.835 $X2=8.47 $Y2=2.95
r207 7 51 400 $w=1.7e-07 $l=4.93559e-07 $layer=licon1_PDIFF $count=1 $X=8.345
+ $Y=1.835 $X2=8.47 $Y2=2.27
r208 6 47 600 $w=1.7e-07 $l=1.00256e-06 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.835 $X2=7.39 $Y2=2.77
r209 5 43 600 $w=1.7e-07 $l=1.01184e-06 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.835 $X2=6.51 $Y2=2.77
r210 4 39 600 $w=1.7e-07 $l=1.05565e-06 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.835 $X2=5.63 $Y2=2.83
r211 3 35 600 $w=1.7e-07 $l=5.17446e-07 $layer=licon1_PDIFF $count=1 $X=4.33
+ $Y=1.795 $X2=4.475 $Y2=2.245
r212 2 31 600 $w=1.7e-07 $l=3.7888e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.795 $X2=1.775 $Y2=2.085
r213 1 27 600 $w=1.7e-07 $l=4.78435e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=2.365 $X2=0.305 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_606_359# 1 2 7 9 14
c33 7 0 9.7377e-20 $X=4.835 $Y=1.86
r34 14 17 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5 $Y=1.86 $X2=5
+ $Y2=2.005
r35 9 12 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=3.18 $Y=1.86 $X2=3.18
+ $Y2=1.95
r36 8 9 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.32 $Y=1.86 $X2=3.18
+ $Y2=1.86
r37 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=1.86 $X2=5
+ $Y2=1.86
r38 7 8 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=4.835 $Y=1.86
+ $X2=3.32 $Y2=1.86
r39 2 17 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.86
+ $Y=1.795 $X2=5 $Y2=2.005
r40 1 12 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.795 $X2=3.155 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%Q 1 2 10 12 13 15 18
c28 13 0 2.67944e-20 $X=6.925 $Y=1.815
c29 12 0 1.4541e-19 $X=6.96 $Y=1.98
r30 15 18 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6.93 $Y=0.925
+ $X2=6.93 $Y2=0.505
r31 12 13 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=1.98
+ $X2=6.925 $Y2=1.815
r32 10 13 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.88 $Y=1.155
+ $X2=6.88 $Y2=1.815
r33 9 15 4.05489 $w=2.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.93 $Y=1.02 $X2=6.93
+ $Y2=0.925
r34 9 10 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.93 $Y=1.02
+ $X2=6.93 $Y2=1.155
r35 2 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.835 $X2=6.96 $Y2=1.98
r36 1 18 91 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=2 $X=6.82
+ $Y=0.3 $X2=6.96 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%Q_N 1 2 7 8 9 10 11 18
r18 11 32 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=8.915 $Y=2.775
+ $X2=8.915 $Y2=2.91
r19 10 11 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=8.915 $Y=2.405
+ $X2=8.915 $Y2=2.775
r20 9 10 20.4078 $w=2.38e-07 $l=4.25e-07 $layer=LI1_cond $X=8.915 $Y=1.98
+ $X2=8.915 $Y2=2.405
r21 8 9 15.1258 $w=2.38e-07 $l=3.15e-07 $layer=LI1_cond $X=8.915 $Y=1.665
+ $X2=8.915 $Y2=1.98
r22 7 8 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=8.915 $Y=1.295
+ $X2=8.915 $Y2=1.665
r23 7 18 42.0162 $w=2.38e-07 $l=8.75e-07 $layer=LI1_cond $X=8.915 $Y=1.295
+ $X2=8.915 $Y2=0.42
r24 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.835 $X2=8.9 $Y2=2.91
r25 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.835 $X2=8.9 $Y2=1.98
r26 1 18 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=8.76
+ $Y=0.27 $X2=8.9 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 46 48
+ 50 52 54 59 64 72 77 82 91 94 97 100 103 107
r112 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r113 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r114 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r115 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r116 94 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r117 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r118 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r119 86 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r120 86 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r121 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r122 83 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=0
+ $X2=8.45 $Y2=0
r123 83 85 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.615 $Y=0
+ $X2=8.88 $Y2=0
r124 82 106 4.38699 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=9.402 $Y2=0
r125 82 85 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r126 81 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r127 81 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r128 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r129 78 100 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.44 $Y2=0
r130 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.92 $Y2=0
r131 77 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=0
+ $X2=8.45 $Y2=0
r132 77 80 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.285 $Y=0
+ $X2=7.92 $Y2=0
r133 76 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r134 76 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r135 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r136 73 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=0 $X2=6.46
+ $Y2=0
r137 73 75 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.625 $Y=0
+ $X2=6.96 $Y2=0
r138 72 100 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.285 $Y=0
+ $X2=7.44 $Y2=0
r139 72 75 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.285 $Y=0
+ $X2=6.96 $Y2=0
r140 71 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r141 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r142 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r143 67 70 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r144 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r145 65 94 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.655
+ $Y2=0
r146 65 67 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=5.04 $Y2=0
r147 64 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.46
+ $Y2=0
r148 64 70 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6
+ $Y2=0
r149 63 95 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r150 63 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r151 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r152 60 91 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.685
+ $Y2=0
r153 60 62 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=2.16 $Y2=0
r154 59 94 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.545 $Y=0 $X2=4.655
+ $Y2=0
r155 59 62 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=4.545 $Y=0
+ $X2=2.16 $Y2=0
r156 58 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r157 58 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r158 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r159 55 88 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r160 55 57 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=1.2
+ $Y2=0
r161 54 91 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.685
+ $Y2=0
r162 54 57 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.2
+ $Y2=0
r163 52 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r164 52 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r165 48 106 3.05085 $w=2.9e-07 $l=1.07912e-07 $layer=LI1_cond $X=9.35 $Y=0.085
+ $X2=9.402 $Y2=0
r166 48 50 13.114 $w=2.88e-07 $l=3.3e-07 $layer=LI1_cond $X=9.35 $Y=0.085
+ $X2=9.35 $Y2=0.415
r167 44 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=0.085
+ $X2=8.45 $Y2=0
r168 44 46 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=8.45 $Y=0.085
+ $X2=8.45 $Y2=0.59
r169 40 42 20.2607 $w=3.08e-07 $l=5.45e-07 $layer=LI1_cond $X=7.44 $Y=0.445
+ $X2=7.44 $Y2=0.99
r170 38 100 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0
r171 38 40 13.3832 $w=3.08e-07 $l=3.6e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0.445
r172 34 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=0.085
+ $X2=6.46 $Y2=0
r173 34 36 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.46 $Y=0.085
+ $X2=6.46 $Y2=0.445
r174 30 94 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0
r175 30 32 26.9776 $w=2.18e-07 $l=5.15e-07 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0.6
r176 26 91 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0
r177 26 28 41.3832 $w=2.18e-07 $l=7.9e-07 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0.875
r178 22 88 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r179 22 24 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.915
r180 7 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.19
+ $Y=0.27 $X2=9.33 $Y2=0.415
r181 6 46 182 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.27 $X2=8.45 $Y2=0.59
r182 5 42 182 $w=1.7e-07 $l=8.05357e-07 $layer=licon1_NDIFF $count=1 $X=7.25
+ $Y=0.3 $X2=7.5 $Y2=0.99
r183 5 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.25
+ $Y=0.3 $X2=7.39 $Y2=0.445
r184 4 36 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.3 $X2=6.46 $Y2=0.445
r185 3 32 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=4.5
+ $Y=0.405 $X2=4.64 $Y2=0.6
r186 2 28 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.72 $X2=1.67 $Y2=0.875
r187 1 24 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.72 $X2=0.275 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_508_155# 1 2 9 11 13
r26 11 13 89.3434 $w=1.78e-07 $l=1.45e-06 $layer=LI1_cond $X=2.76 $Y=0.705
+ $X2=4.21 $Y2=0.705
r27 7 11 6.86909 $w=1.8e-07 $l=1.43091e-07 $layer=LI1_cond $X=2.655 $Y=0.795
+ $X2=2.76 $Y2=0.705
r28 7 9 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=2.655 $Y=0.795
+ $X2=2.655 $Y2=0.985
r29 2 13 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=4.065
+ $Y=0.405 $X2=4.21 $Y2=0.7
r30 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.775 $X2=2.665 $Y2=0.985
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBN_2%A_677_155# 1 2 7 13
r19 11 13 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=5.085 $Y=0.965
+ $X2=5.085 $Y2=0.62
r20 7 11 7.27304 $w=1.9e-07 $l=1.91703e-07 $layer=LI1_cond $X=4.935 $Y=1.06
+ $X2=5.085 $Y2=0.965
r21 7 9 77.6364 $w=1.88e-07 $l=1.33e-06 $layer=LI1_cond $X=4.935 $Y=1.06
+ $X2=3.605 $Y2=1.06
r22 2 13 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.405 $X2=5.07 $Y2=0.62
r23 1 9 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=3.385
+ $Y=0.775 $X2=3.605 $Y2=1.05
.ends

