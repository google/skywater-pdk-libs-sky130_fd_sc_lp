* File: sky130_fd_sc_lp__a41oi_2.spice
* Created: Wed Sep  2 09:29:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41oi_2.pex.spice"
.subckt sky130_fd_sc_lp__a41oi_2  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1011 N_Y_M1011_d N_B1_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_Y_M1011_d N_B1_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_318_69#_M1004_d N_A1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1016 N_A_318_69#_M1016_d N_A1_M1016_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1002 N_A_318_69#_M1016_d N_A2_M1002_g N_A_577_69#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1014 N_A_318_69#_M1014_d N_A2_M1014_g N_A_577_69#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2814 AS=0.1176 PD=2.35 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6
+ SA=75001.5 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1005 N_A_788_69#_M1005_d N_A3_M1005_g N_A_577_69#_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2814 AS=0.1176 PD=2.35 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6
+ SA=75000.3 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1017 N_A_788_69#_M1017_d N_A3_M1017_g N_A_577_69#_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A4_M1009_g N_A_788_69#_M1017_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1009_d N_A4_M1019_g N_A_788_69#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_103_367#_M1001_d N_B1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2 SB=75005
+ A=0.189 P=2.82 MULT=1
MM1007 N_A_103_367#_M1007_d N_B1_M1007_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1000 N_A_103_367#_M1007_d N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.28035 PD=1.54 PS=1.705 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75001.1 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1015 N_A_103_367#_M1015_d N_A1_M1015_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.28035 PD=1.54 PS=1.705 NRD=0 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75003.5 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_A2_M1010_g N_A_103_367#_M1015_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.5418 AS=0.1764 PD=2.12 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75002.1 SB=75003.1 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1010_d N_A2_M1018_g N_A_103_367#_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.5418 AS=0.1764 PD=2.12 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.1
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A3_M1006_g N_A_103_367#_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2835 AS=0.1764 PD=1.71 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75003.5 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1006_d N_A3_M1008_g N_A_103_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2835 AS=0.1764 PD=1.71 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A4_M1003_g N_A_103_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1003_d N_A4_M1013_g N_A_103_367#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__a41oi_2.pxi.spice"
*
.ends
*
*
