* File: sky130_fd_sc_lp__o21a_0.spice
* Created: Fri Aug 28 11:03:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21a_0.pex.spice"
.subckt sky130_fd_sc_lp__o21a_0  VNB VPB B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_80_23#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_300_58#_M1002_d N_B1_M1002_g N_A_80_23#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_300_58#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_300_58#_M1001_d N_A1_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_23#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1072 AS=0.1696 PD=0.975 PS=1.81 NRD=13.8491 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1006 N_A_80_23#_M1006_d N_B1_M1006_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1072 AS=0.1072 PD=0.975 PS=0.975 NRD=0 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1005 A_337_483# N_A2_M1005_g N_A_80_23#_M1006_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1072 PD=0.85 PS=0.975 NRD=15.3857 NRS=16.9223 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_337_483# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__o21a_0.pxi.spice"
*
.ends
*
*
