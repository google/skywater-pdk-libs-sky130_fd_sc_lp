* File: sky130_fd_sc_lp__buf_4.pxi.spice
* Created: Wed Sep  2 09:35:02 2020
* 
x_PM_SKY130_FD_SC_LP__BUF_4%A_122_23# N_A_122_23#_M1001_d N_A_122_23#_M1000_d
+ N_A_122_23#_M1002_g N_A_122_23#_M1004_g N_A_122_23#_M1003_g
+ N_A_122_23#_M1005_g N_A_122_23#_M1006_g N_A_122_23#_M1008_g
+ N_A_122_23#_M1007_g N_A_122_23#_M1009_g N_A_122_23#_c_114_p N_A_122_23#_c_61_n
+ N_A_122_23#_c_62_n N_A_122_23#_c_63_n N_A_122_23#_c_137_p N_A_122_23#_c_72_n
+ N_A_122_23#_c_91_p N_A_122_23#_c_64_n N_A_122_23#_c_73_n N_A_122_23#_c_65_n
+ N_A_122_23#_c_66_n PM_SKY130_FD_SC_LP__BUF_4%A_122_23#
x_PM_SKY130_FD_SC_LP__BUF_4%A N_A_M1001_g N_A_M1000_g A N_A_c_163_n N_A_c_164_n
+ PM_SKY130_FD_SC_LP__BUF_4%A
x_PM_SKY130_FD_SC_LP__BUF_4%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_M1009_d
+ N_VPWR_c_188_n N_VPWR_c_189_n N_VPWR_c_190_n N_VPWR_c_191_n N_VPWR_c_192_n
+ N_VPWR_c_193_n VPWR N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_187_n
+ N_VPWR_c_197_n N_VPWR_c_198_n PM_SKY130_FD_SC_LP__BUF_4%VPWR
x_PM_SKY130_FD_SC_LP__BUF_4%X N_X_M1002_s N_X_M1006_s N_X_M1004_s N_X_M1008_s
+ N_X_c_237_n N_X_c_242_n N_X_c_243_n N_X_c_286_p N_X_c_275_n N_X_c_238_n
+ N_X_c_244_n N_X_c_288_p N_X_c_279_n N_X_c_239_n N_X_c_245_n X X N_X_c_240_n X
+ PM_SKY130_FD_SC_LP__BUF_4%X
x_PM_SKY130_FD_SC_LP__BUF_4%VGND N_VGND_M1002_d N_VGND_M1003_d N_VGND_M1007_d
+ N_VGND_c_293_n N_VGND_c_294_n N_VGND_c_295_n N_VGND_c_296_n N_VGND_c_297_n
+ N_VGND_c_298_n VGND N_VGND_c_299_n N_VGND_c_300_n N_VGND_c_301_n
+ N_VGND_c_302_n N_VGND_c_303_n PM_SKY130_FD_SC_LP__BUF_4%VGND
cc_1 VNB N_A_122_23#_M1002_g 0.0270565f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.665
cc_2 VNB N_A_122_23#_M1003_g 0.0222422f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.665
cc_3 VNB N_A_122_23#_M1006_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=0.665
cc_4 VNB N_A_122_23#_M1007_g 0.0225128f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=0.665
cc_5 VNB N_A_122_23#_c_61_n 0.0023443f $X=-0.19 $Y=-0.245 $X2=2.122 $Y2=1.415
cc_6 VNB N_A_122_23#_c_62_n 4.61888e-19 $X=-0.19 $Y=-0.245 $X2=2.122 $Y2=1.755
cc_7 VNB N_A_122_23#_c_63_n 0.0075508f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=0.945
cc_8 VNB N_A_122_23#_c_64_n 0.0230171f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=0.42
cc_9 VNB N_A_122_23#_c_65_n 0.00146737f $X=-0.19 $Y=-0.245 $X2=2.122 $Y2=1.51
cc_10 VNB N_A_122_23#_c_66_n 0.0663285f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.51
cc_11 VNB N_A_M1000_g 0.00933198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A 0.016977f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.665
cc_13 VNB N_A_c_163_n 0.0369434f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.675
cc_14 VNB N_A_c_164_n 0.023123f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.465
cc_15 VNB N_VPWR_c_187_n 0.123877f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.51
cc_16 VNB N_X_c_237_n 0.00169931f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.465
cc_17 VNB N_X_c_238_n 0.00568171f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=1.675
cc_18 VNB N_X_c_239_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.51
cc_19 VNB N_X_c_240_n 0.0179576f $X=-0.19 $Y=-0.245 $X2=2.122 $Y2=1.605
cc_20 VNB X 0.0246601f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=0.945
cc_21 VNB N_VGND_c_293_n 0.0289266f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.465
cc_22 VNB N_VGND_c_294_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_295_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_296_n 6.09197e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_297_n 0.011849f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=0.665
cc_26 VNB N_VGND_c_298_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=0.665
cc_27 VNB N_VGND_c_299_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.345
cc_28 VNB N_VGND_c_300_n 0.0154417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_301_n 0.176615f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.51
cc_30 VNB N_VGND_c_302_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.51
cc_31 VNB N_VGND_c_303_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.51
cc_32 VPB N_A_122_23#_M1004_g 0.0212719f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.465
cc_33 VPB N_A_122_23#_M1005_g 0.0179927f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.465
cc_34 VPB N_A_122_23#_M1008_g 0.018006f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=2.465
cc_35 VPB N_A_122_23#_M1009_g 0.0178566f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=2.465
cc_36 VPB N_A_122_23#_c_62_n 9.33202e-19 $X=-0.19 $Y=1.655 $X2=2.122 $Y2=1.755
cc_37 VPB N_A_122_23#_c_72_n 0.0136514f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=1.84
cc_38 VPB N_A_122_23#_c_73_n 0.0435297f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=1.98
cc_39 VPB N_A_122_23#_c_66_n 0.0108382f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=1.51
cc_40 VPB N_A_M1000_g 0.0258866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_188_n 0.0399019f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.465
cc_42 VPB N_VPWR_c_189_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.665
cc_43 VPB N_VPWR_c_190_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.465
cc_44 VPB N_VPWR_c_191_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_192_n 0.011849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_193_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=1.345
cc_47 VPB N_VPWR_c_194_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=2.465
cc_48 VPB N_VPWR_c_195_n 0.0153759f $X=-0.19 $Y=1.655 $X2=1.885 $Y2=1.51
cc_49 VPB N_VPWR_c_187_n 0.0527168f $X=-0.19 $Y=1.655 $X2=1.885 $Y2=1.51
cc_50 VPB N_VPWR_c_197_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.122 $Y2=1.415
cc_51 VPB N_VPWR_c_198_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=0.945
cc_52 VPB N_X_c_242_n 0.00169931f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.345
cc_53 VPB N_X_c_243_n 0.0173337f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=0.665
cc_54 VPB N_X_c_244_n 0.00492295f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=2.465
cc_55 VPB N_X_c_245_n 0.00144314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB X 0.00725612f $X=-0.19 $Y=1.655 $X2=2.525 $Y2=0.945
cc_57 N_A_122_23#_M1009_g N_A_M1000_g 0.0230859f $X=1.975 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A_122_23#_c_62_n N_A_M1000_g 0.00339135f $X=2.122 $Y=1.755 $X2=0 $Y2=0
cc_59 N_A_122_23#_c_72_n N_A_M1000_g 0.0158043f $X=2.525 $Y=1.84 $X2=0 $Y2=0
cc_60 N_A_122_23#_M1007_g A 2.96368e-19 $X=1.975 $Y=0.665 $X2=0 $Y2=0
cc_61 N_A_122_23#_c_61_n A 0.0164786f $X=2.122 $Y=1.415 $X2=0 $Y2=0
cc_62 N_A_122_23#_c_63_n A 0.0304116f $X=2.525 $Y=0.945 $X2=0 $Y2=0
cc_63 N_A_122_23#_c_72_n A 0.0271109f $X=2.525 $Y=1.84 $X2=0 $Y2=0
cc_64 N_A_122_23#_c_65_n A 0.0106379f $X=2.122 $Y=1.51 $X2=0 $Y2=0
cc_65 N_A_122_23#_c_63_n N_A_c_163_n 0.00100493f $X=2.525 $Y=0.945 $X2=0 $Y2=0
cc_66 N_A_122_23#_c_72_n N_A_c_163_n 0.00404874f $X=2.525 $Y=1.84 $X2=0 $Y2=0
cc_67 N_A_122_23#_c_65_n N_A_c_163_n 0.00293382f $X=2.122 $Y=1.51 $X2=0 $Y2=0
cc_68 N_A_122_23#_c_66_n N_A_c_163_n 0.0230859f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_69 N_A_122_23#_M1007_g N_A_c_164_n 0.0230859f $X=1.975 $Y=0.665 $X2=0 $Y2=0
cc_70 N_A_122_23#_c_61_n N_A_c_164_n 0.00538545f $X=2.122 $Y=1.415 $X2=0 $Y2=0
cc_71 N_A_122_23#_c_63_n N_A_c_164_n 0.0115732f $X=2.525 $Y=0.945 $X2=0 $Y2=0
cc_72 N_A_122_23#_c_72_n N_VPWR_M1009_d 5.5277e-19 $X=2.525 $Y=1.84 $X2=0 $Y2=0
cc_73 N_A_122_23#_c_91_p N_VPWR_M1009_d 0.00125049f $X=2.22 $Y=1.84 $X2=0 $Y2=0
cc_74 N_A_122_23#_M1004_g N_VPWR_c_188_n 0.0150803f $X=0.685 $Y=2.465 $X2=0
+ $Y2=0
cc_75 N_A_122_23#_M1005_g N_VPWR_c_188_n 7.21513e-19 $X=1.115 $Y=2.465 $X2=0
+ $Y2=0
cc_76 N_A_122_23#_M1004_g N_VPWR_c_189_n 0.00486043f $X=0.685 $Y=2.465 $X2=0
+ $Y2=0
cc_77 N_A_122_23#_M1005_g N_VPWR_c_189_n 0.00486043f $X=1.115 $Y=2.465 $X2=0
+ $Y2=0
cc_78 N_A_122_23#_M1004_g N_VPWR_c_190_n 7.21513e-19 $X=0.685 $Y=2.465 $X2=0
+ $Y2=0
cc_79 N_A_122_23#_M1005_g N_VPWR_c_190_n 0.0140168f $X=1.115 $Y=2.465 $X2=0
+ $Y2=0
cc_80 N_A_122_23#_M1008_g N_VPWR_c_190_n 0.0140168f $X=1.545 $Y=2.465 $X2=0
+ $Y2=0
cc_81 N_A_122_23#_M1009_g N_VPWR_c_190_n 7.21513e-19 $X=1.975 $Y=2.465 $X2=0
+ $Y2=0
cc_82 N_A_122_23#_M1008_g N_VPWR_c_191_n 7.27171e-19 $X=1.545 $Y=2.465 $X2=0
+ $Y2=0
cc_83 N_A_122_23#_M1009_g N_VPWR_c_191_n 0.0141821f $X=1.975 $Y=2.465 $X2=0
+ $Y2=0
cc_84 N_A_122_23#_c_72_n N_VPWR_c_191_n 0.00606161f $X=2.525 $Y=1.84 $X2=0 $Y2=0
cc_85 N_A_122_23#_c_91_p N_VPWR_c_191_n 0.0121776f $X=2.22 $Y=1.84 $X2=0 $Y2=0
cc_86 N_A_122_23#_M1008_g N_VPWR_c_194_n 0.00486043f $X=1.545 $Y=2.465 $X2=0
+ $Y2=0
cc_87 N_A_122_23#_M1009_g N_VPWR_c_194_n 0.00486043f $X=1.975 $Y=2.465 $X2=0
+ $Y2=0
cc_88 N_A_122_23#_c_73_n N_VPWR_c_195_n 0.0178111f $X=2.62 $Y=1.98 $X2=0 $Y2=0
cc_89 N_A_122_23#_M1000_d N_VPWR_c_187_n 0.00371702f $X=2.48 $Y=1.835 $X2=0
+ $Y2=0
cc_90 N_A_122_23#_M1004_g N_VPWR_c_187_n 0.00824727f $X=0.685 $Y=2.465 $X2=0
+ $Y2=0
cc_91 N_A_122_23#_M1005_g N_VPWR_c_187_n 0.00824727f $X=1.115 $Y=2.465 $X2=0
+ $Y2=0
cc_92 N_A_122_23#_M1008_g N_VPWR_c_187_n 0.00824727f $X=1.545 $Y=2.465 $X2=0
+ $Y2=0
cc_93 N_A_122_23#_M1009_g N_VPWR_c_187_n 0.00824727f $X=1.975 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_A_122_23#_c_73_n N_VPWR_c_187_n 0.0100304f $X=2.62 $Y=1.98 $X2=0 $Y2=0
cc_95 N_A_122_23#_M1002_g N_X_c_237_n 0.0169754f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_96 N_A_122_23#_c_114_p N_X_c_237_n 0.00730993f $X=2.025 $Y=1.51 $X2=0 $Y2=0
cc_97 N_A_122_23#_M1004_g N_X_c_242_n 0.0157716f $X=0.685 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_122_23#_c_114_p N_X_c_242_n 0.00730993f $X=2.025 $Y=1.51 $X2=0 $Y2=0
cc_99 N_A_122_23#_M1003_g N_X_c_238_n 0.0141287f $X=1.115 $Y=0.665 $X2=0 $Y2=0
cc_100 N_A_122_23#_M1006_g N_X_c_238_n 0.0137525f $X=1.545 $Y=0.665 $X2=0 $Y2=0
cc_101 N_A_122_23#_M1007_g N_X_c_238_n 0.00131587f $X=1.975 $Y=0.665 $X2=0 $Y2=0
cc_102 N_A_122_23#_c_114_p N_X_c_238_n 0.0625611f $X=2.025 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A_122_23#_c_61_n N_X_c_238_n 0.0133247f $X=2.122 $Y=1.415 $X2=0 $Y2=0
cc_104 N_A_122_23#_c_66_n N_X_c_238_n 0.00497162f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A_122_23#_M1005_g N_X_c_244_n 0.0129249f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_122_23#_M1008_g N_X_c_244_n 0.0128162f $X=1.545 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_122_23#_M1009_g N_X_c_244_n 4.89726e-19 $X=1.975 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_122_23#_c_114_p N_X_c_244_n 0.0625611f $X=2.025 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A_122_23#_c_91_p N_X_c_244_n 0.00911097f $X=2.22 $Y=1.84 $X2=0 $Y2=0
cc_110 N_A_122_23#_c_66_n N_X_c_244_n 0.00497162f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_111 N_A_122_23#_c_114_p N_X_c_239_n 0.0154426f $X=2.025 $Y=1.51 $X2=0 $Y2=0
cc_112 N_A_122_23#_c_66_n N_X_c_239_n 0.00253619f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A_122_23#_c_114_p N_X_c_245_n 0.0154426f $X=2.025 $Y=1.51 $X2=0 $Y2=0
cc_114 N_A_122_23#_c_66_n N_X_c_245_n 0.00253619f $X=1.975 $Y=1.51 $X2=0 $Y2=0
cc_115 N_A_122_23#_M1002_g X 0.0206688f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_116 N_A_122_23#_c_114_p X 0.0147559f $X=2.025 $Y=1.51 $X2=0 $Y2=0
cc_117 N_A_122_23#_c_61_n N_VGND_M1007_d 6.15334e-19 $X=2.122 $Y=1.415 $X2=0
+ $Y2=0
cc_118 N_A_122_23#_c_63_n N_VGND_M1007_d 0.00253014f $X=2.525 $Y=0.945 $X2=0
+ $Y2=0
cc_119 N_A_122_23#_c_137_p N_VGND_M1007_d 0.00123526f $X=2.22 $Y=0.945 $X2=0
+ $Y2=0
cc_120 N_A_122_23#_M1002_g N_VGND_c_293_n 0.0126339f $X=0.685 $Y=0.665 $X2=0
+ $Y2=0
cc_121 N_A_122_23#_M1003_g N_VGND_c_293_n 6.15775e-19 $X=1.115 $Y=0.665 $X2=0
+ $Y2=0
cc_122 N_A_122_23#_M1002_g N_VGND_c_294_n 0.00477554f $X=0.685 $Y=0.665 $X2=0
+ $Y2=0
cc_123 N_A_122_23#_M1003_g N_VGND_c_294_n 0.00477554f $X=1.115 $Y=0.665 $X2=0
+ $Y2=0
cc_124 N_A_122_23#_M1002_g N_VGND_c_295_n 6.15775e-19 $X=0.685 $Y=0.665 $X2=0
+ $Y2=0
cc_125 N_A_122_23#_M1003_g N_VGND_c_295_n 0.0112407f $X=1.115 $Y=0.665 $X2=0
+ $Y2=0
cc_126 N_A_122_23#_M1006_g N_VGND_c_295_n 0.0112407f $X=1.545 $Y=0.665 $X2=0
+ $Y2=0
cc_127 N_A_122_23#_M1007_g N_VGND_c_295_n 6.15775e-19 $X=1.975 $Y=0.665 $X2=0
+ $Y2=0
cc_128 N_A_122_23#_M1006_g N_VGND_c_296_n 5.5495e-19 $X=1.545 $Y=0.665 $X2=0
+ $Y2=0
cc_129 N_A_122_23#_M1007_g N_VGND_c_296_n 0.0100316f $X=1.975 $Y=0.665 $X2=0
+ $Y2=0
cc_130 N_A_122_23#_c_63_n N_VGND_c_296_n 0.00593878f $X=2.525 $Y=0.945 $X2=0
+ $Y2=0
cc_131 N_A_122_23#_c_137_p N_VGND_c_296_n 0.011905f $X=2.22 $Y=0.945 $X2=0 $Y2=0
cc_132 N_A_122_23#_M1006_g N_VGND_c_299_n 0.00477554f $X=1.545 $Y=0.665 $X2=0
+ $Y2=0
cc_133 N_A_122_23#_M1007_g N_VGND_c_299_n 0.00477554f $X=1.975 $Y=0.665 $X2=0
+ $Y2=0
cc_134 N_A_122_23#_c_64_n N_VGND_c_300_n 0.0178111f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_135 N_A_122_23#_M1001_d N_VGND_c_301_n 0.00241995f $X=2.48 $Y=0.245 $X2=0
+ $Y2=0
cc_136 N_A_122_23#_M1002_g N_VGND_c_301_n 0.00825815f $X=0.685 $Y=0.665 $X2=0
+ $Y2=0
cc_137 N_A_122_23#_M1003_g N_VGND_c_301_n 0.00825815f $X=1.115 $Y=0.665 $X2=0
+ $Y2=0
cc_138 N_A_122_23#_M1006_g N_VGND_c_301_n 0.00825815f $X=1.545 $Y=0.665 $X2=0
+ $Y2=0
cc_139 N_A_122_23#_M1007_g N_VGND_c_301_n 0.00825815f $X=1.975 $Y=0.665 $X2=0
+ $Y2=0
cc_140 N_A_122_23#_c_63_n N_VGND_c_301_n 0.00524135f $X=2.525 $Y=0.945 $X2=0
+ $Y2=0
cc_141 N_A_122_23#_c_137_p N_VGND_c_301_n 6.77317e-19 $X=2.22 $Y=0.945 $X2=0
+ $Y2=0
cc_142 N_A_122_23#_c_64_n N_VGND_c_301_n 0.0100304f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_143 N_A_M1000_g N_VPWR_c_191_n 0.0161634f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1000_g N_VPWR_c_195_n 0.00486043f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_VPWR_c_187_n 0.00917987f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_c_164_n N_VGND_c_296_n 0.0116297f $X=2.495 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A_c_164_n N_VGND_c_300_n 0.00477554f $X=2.495 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A_c_164_n N_VGND_c_301_n 0.00552613f $X=2.495 $Y=1.21 $X2=0 $Y2=0
cc_149 N_VPWR_c_187_n N_X_M1004_s 0.00536646f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_150 N_VPWR_c_187_n N_X_M1008_s 0.00536646f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_151 N_VPWR_M1004_d N_X_c_242_n 4.46468e-19 $X=0.325 $Y=1.835 $X2=0 $Y2=0
cc_152 N_VPWR_c_188_n N_X_c_242_n 0.00524802f $X=0.47 $Y=2.2 $X2=0 $Y2=0
cc_153 N_VPWR_M1004_d N_X_c_243_n 0.00268655f $X=0.325 $Y=1.835 $X2=0 $Y2=0
cc_154 N_VPWR_c_188_n N_X_c_243_n 0.0184602f $X=0.47 $Y=2.2 $X2=0 $Y2=0
cc_155 N_VPWR_c_189_n N_X_c_275_n 0.0124525f $X=1.165 $Y=3.33 $X2=0 $Y2=0
cc_156 N_VPWR_c_187_n N_X_c_275_n 0.00730901f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_M1005_d N_X_c_244_n 0.00176461f $X=1.19 $Y=1.835 $X2=0 $Y2=0
cc_158 N_VPWR_c_190_n N_X_c_244_n 0.0170777f $X=1.33 $Y=2.2 $X2=0 $Y2=0
cc_159 N_VPWR_c_194_n N_X_c_279_n 0.0124525f $X=2.025 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_187_n N_X_c_279_n 0.00730901f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_161 N_X_c_237_n N_VGND_M1002_d 4.46468e-19 $X=0.805 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_162 N_X_c_240_n N_VGND_M1002_d 0.00187298f $X=0.302 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_163 N_X_c_238_n N_VGND_M1003_d 0.00176461f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_164 N_X_c_237_n N_VGND_c_293_n 0.00524802f $X=0.805 $Y=1.16 $X2=0 $Y2=0
cc_165 N_X_c_240_n N_VGND_c_293_n 0.0185309f $X=0.302 $Y=1.245 $X2=0 $Y2=0
cc_166 N_X_c_286_p N_VGND_c_294_n 0.0124525f $X=0.9 $Y=0.42 $X2=0 $Y2=0
cc_167 N_X_c_238_n N_VGND_c_295_n 0.0170777f $X=1.665 $Y=1.16 $X2=0 $Y2=0
cc_168 N_X_c_288_p N_VGND_c_299_n 0.0124525f $X=1.76 $Y=0.42 $X2=0 $Y2=0
cc_169 N_X_M1002_s N_VGND_c_301_n 0.00536646f $X=0.76 $Y=0.245 $X2=0 $Y2=0
cc_170 N_X_M1006_s N_VGND_c_301_n 0.00536646f $X=1.62 $Y=0.245 $X2=0 $Y2=0
cc_171 N_X_c_286_p N_VGND_c_301_n 0.00730901f $X=0.9 $Y=0.42 $X2=0 $Y2=0
cc_172 N_X_c_288_p N_VGND_c_301_n 0.00730901f $X=1.76 $Y=0.42 $X2=0 $Y2=0
