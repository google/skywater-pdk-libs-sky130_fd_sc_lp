* File: sky130_fd_sc_lp__nor2_lp2.pxi.spice
* Created: Fri Aug 28 10:53:57 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_LP2%A N_A_M1005_g N_A_M1000_g N_A_c_39_n N_A_M1002_g
+ A A N_A_c_42_n PM_SKY130_FD_SC_LP__NOR2_LP2%A
x_PM_SKY130_FD_SC_LP__NOR2_LP2%B N_B_c_77_n N_B_M1004_g N_B_c_70_n N_B_c_71_n
+ N_B_M1003_g N_B_c_73_n N_B_M1001_g N_B_c_81_n B B B B B N_B_c_76_n
+ PM_SKY130_FD_SC_LP__NOR2_LP2%B
x_PM_SKY130_FD_SC_LP__NOR2_LP2%VPWR N_VPWR_M1005_s N_VPWR_c_112_n N_VPWR_c_113_n
+ VPWR N_VPWR_c_114_n N_VPWR_c_111_n PM_SKY130_FD_SC_LP__NOR2_LP2%VPWR
x_PM_SKY130_FD_SC_LP__NOR2_LP2%Y N_Y_M1002_d N_Y_M1004_d Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__NOR2_LP2%Y
x_PM_SKY130_FD_SC_LP__NOR2_LP2%VGND N_VGND_M1000_s N_VGND_M1001_d N_VGND_c_152_n
+ N_VGND_c_153_n N_VGND_c_154_n N_VGND_c_155_n VGND N_VGND_c_156_n
+ N_VGND_c_157_n PM_SKY130_FD_SC_LP__NOR2_LP2%VGND
cc_1 VNB N_A_M1005_g 0.0111307f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.37
cc_2 VNB N_A_M1000_g 0.0274458f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.77
cc_3 VNB N_A_c_39_n 0.0210976f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=1.255
cc_4 VNB N_A_M1002_g 0.0192706f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.77
cc_5 VNB A 0.0260936f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A_c_42_n 0.0331952f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.255
cc_7 VNB N_B_c_70_n 0.00558371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_71_n 0.00626936f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.18
cc_9 VNB N_B_M1003_g 0.0431429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_73_n 0.00208163f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.255
cc_11 VNB N_B_M1001_g 0.0274385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB B 0.0364239f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_B_c_76_n 0.0430983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_111_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB Y 0.00493081f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.77
cc_16 VNB N_VGND_c_152_n 0.0147687f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.77
cc_17 VNB N_VGND_c_153_n 0.0452411f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=1.255
cc_18 VNB N_VGND_c_154_n 0.0160446f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.18
cc_19 VNB N_VGND_c_155_n 0.0452369f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.77
cc_20 VNB N_VGND_c_156_n 0.0391487f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_21 VNB N_VGND_c_157_n 0.188418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A_M1005_g 0.0326912f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.37
cc_23 VPB A 0.0157628f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_24 VPB N_B_c_77_n 0.0237243f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.51
cc_25 VPB N_B_c_70_n 0.0081775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_B_c_71_n 0.00608227f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.18
cc_27 VPB N_B_c_73_n 0.0128244f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.255
cc_28 VPB N_B_c_81_n 0.00854124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB B 0.0918786f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_30 VPB N_B_c_76_n 0.010505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_112_n 0.0121909f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_113_n 0.0517326f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.77
cc_33 VPB N_VPWR_c_114_n 0.057246f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_34 VPB N_VPWR_c_111_n 0.0778636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB Y 0.0035782f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.77
cc_36 N_A_M1005_g N_B_c_71_n 0.0862721f $X=0.545 $Y=2.37 $X2=0 $Y2=0
cc_37 N_A_c_39_n N_B_c_71_n 0.00878864f $X=0.89 $Y=1.255 $X2=0 $Y2=0
cc_38 A N_B_c_71_n 0.00119296f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_39 N_A_M1002_g N_B_M1003_g 0.0230493f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_40 A N_B_M1003_g 8.96801e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_41 N_A_c_42_n N_B_M1003_g 0.00359846f $X=0.495 $Y=1.255 $X2=0 $Y2=0
cc_42 N_A_M1005_g N_VPWR_c_113_n 0.0239392f $X=0.545 $Y=2.37 $X2=0 $Y2=0
cc_43 A N_VPWR_c_113_n 0.0232372f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_44 N_A_c_42_n N_VPWR_c_113_n 3.28173e-19 $X=0.495 $Y=1.255 $X2=0 $Y2=0
cc_45 N_A_M1005_g N_VPWR_c_114_n 0.00769487f $X=0.545 $Y=2.37 $X2=0 $Y2=0
cc_46 N_A_M1005_g N_VPWR_c_111_n 0.00779694f $X=0.545 $Y=2.37 $X2=0 $Y2=0
cc_47 N_A_M1005_g Y 0.0039042f $X=0.545 $Y=2.37 $X2=0 $Y2=0
cc_48 N_A_M1000_g Y 0.0024689f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_49 N_A_c_39_n Y 0.00461791f $X=0.89 $Y=1.255 $X2=0 $Y2=0
cc_50 N_A_M1002_g Y 0.0168258f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_51 A Y 0.0496026f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_A_c_42_n Y 9.66061e-19 $X=0.495 $Y=1.255 $X2=0 $Y2=0
cc_53 N_A_M1000_g N_VGND_c_153_n 0.0140139f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_54 N_A_M1002_g N_VGND_c_153_n 0.00163467f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_55 A N_VGND_c_153_n 0.0280767f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_c_42_n N_VGND_c_153_n 0.0044847f $X=0.495 $Y=1.255 $X2=0 $Y2=0
cc_57 N_A_M1000_g N_VGND_c_156_n 0.00375057f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_58 N_A_M1002_g N_VGND_c_156_n 0.0043233f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_59 N_A_M1000_g N_VGND_c_157_n 0.00409726f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_VGND_c_157_n 0.00487769f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_61 N_B_c_77_n N_VPWR_c_113_n 0.0027832f $X=1.005 $Y=1.795 $X2=0 $Y2=0
cc_62 N_B_c_77_n N_VPWR_c_114_n 0.00751315f $X=1.005 $Y=1.795 $X2=0 $Y2=0
cc_63 B N_VPWR_c_114_n 0.0231512f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_64 N_B_c_77_n N_VPWR_c_111_n 0.00862493f $X=1.005 $Y=1.795 $X2=0 $Y2=0
cc_65 B N_VPWR_c_111_n 0.0246855f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_66 N_B_c_77_n Y 0.0320519f $X=1.005 $Y=1.795 $X2=0 $Y2=0
cc_67 N_B_c_70_n Y 0.0117133f $X=1.32 $Y=1.72 $X2=0 $Y2=0
cc_68 N_B_c_71_n Y 0.00554503f $X=1.13 $Y=1.72 $X2=0 $Y2=0
cc_69 N_B_M1003_g Y 0.0325474f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_70 N_B_M1001_g Y 0.00269839f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_71 N_B_c_81_n Y 0.00503179f $X=1.395 $Y=1.72 $X2=0 $Y2=0
cc_72 B Y 0.147769f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_73 N_B_c_76_n Y 4.03018e-19 $X=1.875 $Y=1.345 $X2=0 $Y2=0
cc_74 N_B_M1003_g N_VGND_c_155_n 0.00159468f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_75 N_B_M1001_g N_VGND_c_155_n 0.01352f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_76 B N_VGND_c_155_n 0.028459f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_77 N_B_c_76_n N_VGND_c_155_n 0.00141406f $X=1.875 $Y=1.345 $X2=0 $Y2=0
cc_78 N_B_M1003_g N_VGND_c_156_n 0.00392868f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_79 N_B_M1001_g N_VGND_c_156_n 0.00375057f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_80 N_B_M1003_g N_VGND_c_157_n 0.00487769f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_81 N_B_M1001_g N_VGND_c_157_n 0.00409726f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_82 N_VPWR_c_113_n Y 0.0254753f $X=0.28 $Y=2.065 $X2=0 $Y2=0
cc_83 N_VPWR_c_114_n Y 0.0120584f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_84 N_VPWR_c_111_n Y 0.0130683f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_85 Y N_VGND_c_153_n 0.0179348f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_86 Y N_VGND_c_155_n 0.019674f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_87 Y N_VGND_c_156_n 0.0121008f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_88 Y N_VGND_c_157_n 0.0130839f $X=1.115 $Y=0.47 $X2=0 $Y2=0
