* File: sky130_fd_sc_lp__a21oi_0.pex.spice
* Created: Wed Sep  2 09:20:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21OI_0%A2 2 5 7 9 13 16 19 21 22 23 28
c45 21 0 7.11268e-21 $X=0.24 $Y=0.925
r46 22 23 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.665
r47 21 22 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=1.295
r48 21 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r49 17 19 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.36 $Y=2.11
+ $X2=0.565 $Y2=2.11
r50 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r51 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r52 11 28 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.27 $Y=0.915 $X2=0.27
+ $Y2=1.005
r53 11 13 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.27 $Y=0.84
+ $X2=0.605 $Y2=0.84
r54 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.605 $Y=0.765
+ $X2=0.605 $Y2=0.84
r55 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.605 $Y=0.765
+ $X2=0.605 $Y2=0.445
r56 3 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=2.185
+ $X2=0.565 $Y2=2.11
r57 3 5 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.565 $Y=2.185 $X2=0.565
+ $Y2=2.685
r58 2 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.035
+ $X2=0.36 $Y2=2.11
r59 2 16 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=0.36 $Y=2.035
+ $X2=0.36 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_0%A1 2 5 9 11 12 13 14 15 22 31
c49 9 0 3.44349e-20 $X=0.995 $Y=2.685
r50 29 31 0.259705 $w=3.53e-07 $l=8e-09 $layer=LI1_cond $X=0.747 $Y=0.917
+ $X2=0.747 $Y2=0.925
r51 22 24 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.872 $Y=1.32
+ $X2=0.872 $Y2=1.155
r52 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.32 $X2=0.84 $Y2=1.32
r53 15 23 11.1998 $w=3.53e-07 $l=3.45e-07 $layer=LI1_cond $X=0.747 $Y=1.665
+ $X2=0.747 $Y2=1.32
r54 14 23 0.81158 $w=3.53e-07 $l=2.5e-08 $layer=LI1_cond $X=0.747 $Y=1.295
+ $X2=0.747 $Y2=1.32
r55 13 29 1.26606 $w=3.53e-07 $l=3.9e-08 $layer=LI1_cond $X=0.747 $Y=0.878
+ $X2=0.747 $Y2=0.917
r56 13 40 4.78995 $w=3.53e-07 $l=1.38e-07 $layer=LI1_cond $X=0.747 $Y=0.878
+ $X2=0.747 $Y2=0.74
r57 13 14 10.7778 $w=3.53e-07 $l=3.32e-07 $layer=LI1_cond $X=0.747 $Y=0.963
+ $X2=0.747 $Y2=1.295
r58 13 31 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=0.747 $Y=0.963
+ $X2=0.747 $Y2=0.925
r59 12 40 7.10673 $w=2.98e-07 $l=1.85e-07 $layer=LI1_cond $X=0.775 $Y=0.555
+ $X2=0.775 $Y2=0.74
r60 9 11 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.995 $Y=2.685
+ $X2=0.995 $Y2=1.825
r61 5 24 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.995 $Y=0.445
+ $X2=0.995 $Y2=1.155
r62 2 11 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.872 $Y=1.628
+ $X2=0.872 $Y2=1.825
r63 1 22 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.872 $Y=1.352
+ $X2=0.872 $Y2=1.32
r64 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.872 $Y=1.352
+ $X2=0.872 $Y2=1.628
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_0%B1 3 7 9 10 16
r28 13 16 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.425 $Y=1.27
+ $X2=1.62 $Y2=1.27
r29 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.27 $X2=1.62 $Y2=1.27
r30 9 10 10.6025 $w=3.73e-07 $l=3.45e-07 $layer=LI1_cond $X=1.642 $Y=0.925
+ $X2=1.642 $Y2=1.27
r31 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.435
+ $X2=1.425 $Y2=1.27
r32 5 7 640.957 $w=1.5e-07 $l=1.25e-06 $layer=POLY_cond $X=1.425 $Y=1.435
+ $X2=1.425 $Y2=2.685
r33 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.105
+ $X2=1.425 $Y2=1.27
r34 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.425 $Y=1.105
+ $X2=1.425 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_0%A_45_473# 1 2 9 11 12 15
c28 9 0 2.73222e-20 $X=0.35 $Y=2.51
r29 13 15 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=1.212 $Y=2.175
+ $X2=1.212 $Y2=2.51
r30 11 13 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.085 $Y=2.09
+ $X2=1.212 $Y2=2.175
r31 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.085 $Y=2.09
+ $X2=0.475 $Y2=2.09
r32 7 12 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.33 $Y=2.175
+ $X2=0.475 $Y2=2.09
r33 7 9 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=0.33 $Y=2.175
+ $X2=0.33 $Y2=2.51
r34 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=2.365 $X2=1.21 $Y2=2.51
r35 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.365 $X2=0.35 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_0%VPWR 1 8 10 14 15 18
r22 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r24 12 18 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=0.78 $Y2=3.33
r25 12 14 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 10 15 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 10 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 6 18 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r29 6 8 31.3721 $w=2.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.51
r30 1 8 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.64
+ $Y=2.365 $X2=0.78 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_0%Y 1 2 8 9 10 12 15 16 17 18
r30 18 31 9.39684 $w=3.23e-07 $l=2.65e-07 $layer=LI1_cond $X=1.672 $Y=2.775
+ $X2=1.672 $Y2=2.51
r31 17 31 3.72328 $w=3.23e-07 $l=1.05e-07 $layer=LI1_cond $X=1.672 $Y=2.405
+ $X2=1.672 $Y2=2.51
r32 16 17 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.672 $Y=2.035
+ $X2=1.672 $Y2=2.405
r33 15 16 8.29721 $w=4.93e-07 $l=2.85e-07 $layer=LI1_cond $X=1.672 $Y=1.75
+ $X2=1.672 $Y2=2.035
r34 12 14 8.37256 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.217 $Y=0.445
+ $X2=1.217 $Y2=0.61
r35 9 15 4.76901 $w=1.85e-07 $l=1.62e-07 $layer=LI1_cond $X=1.51 $Y=1.657
+ $X2=1.672 $Y2=1.657
r36 9 10 13.4889 $w=1.83e-07 $l=2.25e-07 $layer=LI1_cond $X=1.51 $Y=1.657
+ $X2=1.285 $Y2=1.657
r37 8 10 6.81807 $w=1.85e-07 $l=1.33285e-07 $layer=LI1_cond $X=1.19 $Y=1.565
+ $X2=1.285 $Y2=1.657
r38 8 14 55.7464 $w=1.88e-07 $l=9.55e-07 $layer=LI1_cond $X=1.19 $Y=1.565
+ $X2=1.19 $Y2=0.61
r39 2 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.365 $X2=1.64 $Y2=2.51
r40 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.21 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_0%VGND 1 2 7 9 11 13 15 17 27
r32 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r33 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r34 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r35 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r36 18 23 3.915 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r37 18 20 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=1.2
+ $Y2=0
r38 17 26 4.40486 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.715
+ $Y2=0
r39 17 20 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.2
+ $Y2=0
r40 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r41 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r42 11 26 3.07266 $w=2.95e-07 $l=1.1025e-07 $layer=LI1_cond $X=1.657 $Y=0.085
+ $X2=1.715 $Y2=0
r43 11 13 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=1.657 $Y=0.085
+ $X2=1.657 $Y2=0.445
r44 7 23 3.22816 $w=2.5e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.227 $Y2=0
r45 7 9 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=0.33 $Y=0.085 $X2=0.33
+ $Y2=0.445
r46 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.235 $X2=1.64 $Y2=0.445
r47 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.445
.ends

