* File: sky130_fd_sc_lp__o2bb2ai_4.pxi.spice
* Created: Fri Aug 28 11:12:58 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%B1 N_B1_M1017_g N_B1_M1009_g N_B1_M1019_g
+ N_B1_M1012_g N_B1_M1034_g N_B1_M1036_g N_B1_M1039_g N_B1_M1038_g N_B1_c_166_n
+ N_B1_c_187_p B1 B1 B1 B1 B1 B1 N_B1_c_167_n N_B1_c_168_n N_B1_c_175_n
+ N_B1_c_179_p PM_SKY130_FD_SC_LP__O2BB2AI_4%B1
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%B2 N_B2_M1010_g N_B2_M1005_g N_B2_M1015_g
+ N_B2_M1021_g N_B2_M1029_g N_B2_M1032_g N_B2_M1030_g N_B2_M1037_g B2 B2 B2 B2
+ N_B2_c_290_n PM_SKY130_FD_SC_LP__O2BB2AI_4%B2
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%A_804_39# N_A_804_39#_M1001_s
+ N_A_804_39#_M1018_s N_A_804_39#_M1000_s N_A_804_39#_M1022_s
+ N_A_804_39#_M1007_d N_A_804_39#_M1028_d N_A_804_39#_M1011_g
+ N_A_804_39#_M1002_g N_A_804_39#_M1008_g N_A_804_39#_M1023_g
+ N_A_804_39#_M1013_g N_A_804_39#_M1027_g N_A_804_39#_M1025_g
+ N_A_804_39#_M1031_g N_A_804_39#_c_372_n N_A_804_39#_c_373_n
+ N_A_804_39#_c_383_n N_A_804_39#_c_384_n N_A_804_39#_c_478_p
+ N_A_804_39#_c_385_n N_A_804_39#_c_481_p N_A_804_39#_c_386_n
+ N_A_804_39#_c_482_p N_A_804_39#_c_387_n N_A_804_39#_c_424_p
+ N_A_804_39#_c_483_p N_A_804_39#_c_388_n N_A_804_39#_c_374_n
+ N_A_804_39#_c_375_n N_A_804_39#_c_390_n N_A_804_39#_c_391_n
+ N_A_804_39#_c_422_p N_A_804_39#_c_392_n N_A_804_39#_c_376_n
+ N_A_804_39#_c_393_n N_A_804_39#_c_377_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_4%A_804_39#
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%A1_N N_A1_N_M1000_g N_A1_N_M1003_g
+ N_A1_N_M1006_g N_A1_N_M1004_g N_A1_N_M1022_g N_A1_N_M1024_g N_A1_N_M1026_g
+ N_A1_N_M1035_g N_A1_N_c_562_n A1_N A1_N N_A1_N_c_563_n N_A1_N_c_564_n
+ N_A1_N_c_565_n PM_SKY130_FD_SC_LP__O2BB2AI_4%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%A2_N N_A2_N_c_658_n N_A2_N_M1007_g
+ N_A2_N_M1001_g N_A2_N_c_659_n N_A2_N_M1014_g N_A2_N_M1016_g N_A2_N_c_660_n
+ N_A2_N_M1028_g N_A2_N_M1018_g N_A2_N_c_661_n N_A2_N_M1033_g N_A2_N_M1020_g
+ N_A2_N_c_654_n A2_N A2_N N_A2_N_c_655_n N_A2_N_c_656_n N_A2_N_c_657_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_4%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%VPWR N_VPWR_M1009_d N_VPWR_M1012_d
+ N_VPWR_M1038_d N_VPWR_M1008_s N_VPWR_M1025_s N_VPWR_M1006_d N_VPWR_M1026_d
+ N_VPWR_M1014_s N_VPWR_M1033_s N_VPWR_c_736_n N_VPWR_c_737_n N_VPWR_c_738_n
+ N_VPWR_c_739_n N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_742_n N_VPWR_c_743_n
+ N_VPWR_c_744_n N_VPWR_c_745_n N_VPWR_c_746_n N_VPWR_c_747_n N_VPWR_c_748_n
+ N_VPWR_c_749_n N_VPWR_c_750_n N_VPWR_c_751_n N_VPWR_c_752_n VPWR
+ N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_755_n N_VPWR_c_756_n N_VPWR_c_757_n
+ N_VPWR_c_758_n N_VPWR_c_759_n N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_735_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%A_132_367# N_A_132_367#_M1009_s
+ N_A_132_367#_M1036_s N_A_132_367#_M1021_s N_A_132_367#_M1037_s
+ N_A_132_367#_c_895_n N_A_132_367#_c_922_n N_A_132_367#_c_905_n
+ N_A_132_367#_c_910_n N_A_132_367#_c_927_n N_A_132_367#_c_911_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_4%A_132_367#
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%Y N_Y_M1011_s N_Y_M1027_s N_Y_M1005_d
+ N_Y_M1032_d N_Y_M1002_d N_Y_M1013_d N_Y_c_936_n N_Y_c_964_n N_Y_c_965_n
+ N_Y_c_993_n N_Y_c_940_n N_Y_c_937_n N_Y_c_997_n N_Y_c_979_n N_Y_c_938_n
+ N_Y_c_941_n Y Y Y Y Y PM_SKY130_FD_SC_LP__O2BB2AI_4%Y
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%A_35_65# N_A_35_65#_M1017_d N_A_35_65#_M1019_d
+ N_A_35_65#_M1010_d N_A_35_65#_M1029_d N_A_35_65#_M1039_d N_A_35_65#_M1023_d
+ N_A_35_65#_M1031_d N_A_35_65#_c_1021_n N_A_35_65#_c_1022_n N_A_35_65#_c_1023_n
+ N_A_35_65#_c_1024_n N_A_35_65#_c_1025_n N_A_35_65#_c_1026_n
+ N_A_35_65#_c_1027_n N_A_35_65#_c_1028_n N_A_35_65#_c_1029_n
+ N_A_35_65#_c_1052_n N_A_35_65#_c_1053_n N_A_35_65#_c_1030_n
+ N_A_35_65#_c_1031_n N_A_35_65#_c_1080_n N_A_35_65#_c_1032_n
+ N_A_35_65#_c_1033_n N_A_35_65#_c_1034_n N_A_35_65#_c_1035_n
+ N_A_35_65#_c_1036_n N_A_35_65#_c_1057_n N_A_35_65#_c_1037_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_4%A_35_65#
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%VGND N_VGND_M1017_s N_VGND_M1034_s
+ N_VGND_M1015_s N_VGND_M1030_s N_VGND_M1003_s N_VGND_M1024_s N_VGND_c_1138_n
+ N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n
+ N_VGND_c_1143_n N_VGND_c_1144_n N_VGND_c_1145_n N_VGND_c_1146_n
+ N_VGND_c_1147_n N_VGND_c_1148_n N_VGND_c_1149_n N_VGND_c_1150_n
+ N_VGND_c_1151_n N_VGND_c_1152_n VGND N_VGND_c_1153_n N_VGND_c_1154_n
+ N_VGND_c_1155_n N_VGND_c_1156_n N_VGND_c_1157_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_4%VGND
x_PM_SKY130_FD_SC_LP__O2BB2AI_4%A_1235_65# N_A_1235_65#_M1003_d
+ N_A_1235_65#_M1004_d N_A_1235_65#_M1035_d N_A_1235_65#_M1016_d
+ N_A_1235_65#_M1020_d N_A_1235_65#_c_1273_n N_A_1235_65#_c_1274_n
+ N_A_1235_65#_c_1299_n N_A_1235_65#_c_1275_n N_A_1235_65#_c_1276_n
+ N_A_1235_65#_c_1277_n N_A_1235_65#_c_1278_n N_A_1235_65#_c_1279_n
+ N_A_1235_65#_c_1280_n N_A_1235_65#_c_1281_n N_A_1235_65#_c_1282_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_4%A_1235_65#
cc_1 VNB N_B1_M1017_g 0.0259913f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.745
cc_2 VNB N_B1_M1019_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.745
cc_3 VNB N_B1_M1034_g 0.0192613f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=0.745
cc_4 VNB N_B1_M1039_g 0.0184588f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=0.745
cc_5 VNB N_B1_c_166_n 0.00887859f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.535
cc_6 VNB N_B1_c_167_n 0.0607522f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.51
cc_7 VNB N_B1_c_168_n 0.0290123f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.51
cc_8 VNB N_B2_M1010_g 0.0192613f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.745
cc_9 VNB N_B2_M1015_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.745
cc_10 VNB N_B2_M1029_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=0.745
cc_11 VNB N_B2_M1030_g 0.0200792f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=0.745
cc_12 VNB B2 0.00263794f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.51
cc_13 VNB N_B2_c_290_n 0.0697334f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.51
cc_14 VNB N_A_804_39#_M1011_g 0.0194898f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.675
cc_15 VNB N_A_804_39#_M1023_g 0.0203562f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.535
cc_16 VNB N_A_804_39#_M1027_g 0.0210569f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.51
cc_17 VNB N_A_804_39#_M1031_g 0.0251932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_804_39#_c_372_n 0.0015582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_804_39#_c_373_n 6.64882e-19 $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.51
cc_20 VNB N_A_804_39#_c_374_n 0.0111862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_804_39#_c_375_n 0.0197325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_804_39#_c_376_n 0.00228483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_804_39#_c_377_n 0.0784593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_N_M1003_g 0.0248286f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_25 VNB N_A1_N_M1004_g 0.0198186f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.465
cc_26 VNB N_A1_N_M1024_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=2.465
cc_27 VNB N_A1_N_M1035_g 0.0194899f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_28 VNB N_A1_N_c_562_n 0.00136137f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.645
cc_29 VNB N_A1_N_c_563_n 0.089903f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.51
cc_30 VNB N_A1_N_c_564_n 0.0150191f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.51
cc_31 VNB N_A1_N_c_565_n 6.2384e-19 $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.51
cc_32 VNB N_A2_N_M1001_g 0.0194885f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_33 VNB N_A2_N_M1016_g 0.0184296f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.675
cc_34 VNB N_A2_N_M1018_g 0.0194148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_N_M1020_g 0.0234315f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=0.745
cc_36 VNB N_A2_N_c_654_n 0.00160869f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_37 VNB N_A2_N_c_655_n 0.0723605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A2_N_c_656_n 0.00280418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A2_N_c_657_n 0.00342799f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.51
cc_40 VNB N_VPWR_c_735_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_936_n 0.00326045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_937_n 0.00554228f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.51
cc_43 VNB N_Y_c_938_n 0.00342442f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.95
cc_44 VNB N_A_35_65#_c_1021_n 0.0310467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_35_65#_c_1022_n 0.00313953f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=0.745
cc_46 VNB N_A_35_65#_c_1023_n 0.0150832f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=0.745
cc_47 VNB N_A_35_65#_c_1024_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=2.465
cc_48 VNB N_A_35_65#_c_1025_n 0.00529219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_35_65#_c_1026_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.51
cc_50 VNB N_A_35_65#_c_1027_n 0.0030484f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.645
cc_51 VNB N_A_35_65#_c_1028_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_52 VNB N_A_35_65#_c_1029_n 0.0106316f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.95
cc_53 VNB N_A_35_65#_c_1030_n 0.00281114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_35_65#_c_1031_n 0.00225111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_35_65#_c_1032_n 0.00675882f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.51
cc_56 VNB N_A_35_65#_c_1033_n 0.00572422f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.51
cc_57 VNB N_A_35_65#_c_1034_n 0.00143873f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.51
cc_58 VNB N_A_35_65#_c_1035_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_35_65#_c_1036_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.51
cc_60 VNB N_A_35_65#_c_1037_n 0.00224938f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.51
cc_61 VNB N_VGND_c_1138_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.675
cc_62 VNB N_VGND_c_1139_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=3.605 $Y2=1.295
cc_63 VNB N_VGND_c_1140_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=1.675
cc_64 VNB N_VGND_c_1141_n 0.00457468f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.535
cc_65 VNB N_VGND_c_1142_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1143_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.535
cc_67 VNB N_VGND_c_1144_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.95
cc_68 VNB N_VGND_c_1145_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.95
cc_69 VNB N_VGND_c_1146_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.95
cc_70 VNB N_VGND_c_1147_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1148_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1149_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1150_n 0.00600906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1151_n 0.0741762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1152_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1153_n 0.0175526f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.51
cc_77 VNB N_VGND_c_1154_n 0.0566869f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.51
cc_78 VNB N_VGND_c_1155_n 0.530919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1156_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1157_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1235_65#_c_1273_n 0.00180138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1235_65#_c_1274_n 0.00732566f $X=-0.19 $Y=-0.245 $X2=1.375
+ $Y2=0.745
cc_83 VNB N_A_1235_65#_c_1275_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1235_65#_c_1276_n 0.00654355f $X=-0.19 $Y=-0.245 $X2=3.605
+ $Y2=0.745
cc_85 VNB N_A_1235_65#_c_1277_n 0.00257379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1235_65#_c_1278_n 0.00185825f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=1.535
cc_87 VNB N_A_1235_65#_c_1279_n 0.0128308f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.535
cc_88 VNB N_A_1235_65#_c_1280_n 0.0185206f $X=-0.19 $Y=-0.245 $X2=1.235
+ $Y2=1.645
cc_89 VNB N_A_1235_65#_c_1281_n 0.0024549f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_90 VNB N_A_1235_65#_c_1282_n 0.00181463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VPB N_B1_M1009_g 0.0255701f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_92 VPB N_B1_M1012_g 0.017861f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.465
cc_93 VPB N_B1_M1036_g 0.0184774f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=2.465
cc_94 VPB N_B1_M1038_g 0.0179515f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=2.465
cc_95 VPB N_B1_c_167_n 0.0128777f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=1.51
cc_96 VPB N_B1_c_168_n 0.00645128f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=1.51
cc_97 VPB N_B1_c_175_n 0.00236492f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=1.51
cc_98 VPB N_B2_M1005_g 0.0183737f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_99 VPB N_B2_M1021_g 0.017887f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.465
cc_100 VPB N_B2_M1032_g 0.0178862f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=2.465
cc_101 VPB N_B2_M1037_g 0.0186048f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=2.465
cc_102 VPB B2 0.0107514f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.51
cc_103 VPB N_B2_c_290_n 0.0152268f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.51
cc_104 VPB N_A_804_39#_M1002_g 0.018045f $X=-0.19 $Y=1.655 $X2=3.605 $Y2=1.295
cc_105 VPB N_A_804_39#_M1008_g 0.0180054f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=1.675
cc_106 VPB N_A_804_39#_M1013_g 0.0180101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_804_39#_M1025_g 0.0214351f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.95
cc_108 VPB N_A_804_39#_c_373_n 0.00204767f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.51
cc_109 VPB N_A_804_39#_c_383_n 0.00832911f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.51
cc_110 VPB N_A_804_39#_c_384_n 5.30069e-19 $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.51
cc_111 VPB N_A_804_39#_c_385_n 0.0030484f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=1.295
cc_112 VPB N_A_804_39#_c_386_n 0.00748889f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=2.04
cc_113 VPB N_A_804_39#_c_387_n 0.00313447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_804_39#_c_388_n 0.0161202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_804_39#_c_375_n 0.00558299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_804_39#_c_390_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_804_39#_c_391_n 0.00143549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_804_39#_c_392_n 0.00143553f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_804_39#_c_393_n 0.00134162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_804_39#_c_377_n 0.0183819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A1_N_M1000_g 0.0207909f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.745
cc_122 VPB N_A1_N_M1006_g 0.0179297f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=0.745
cc_123 VPB N_A1_N_M1022_g 0.0179297f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=0.745
cc_124 VPB N_A1_N_M1026_g 0.0208607f $X=-0.19 $Y=1.655 $X2=3.605 $Y2=0.745
cc_125 VPB N_A1_N_c_563_n 0.0220624f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.51
cc_126 VPB N_A2_N_c_658_n 0.0177076f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.345
cc_127 VPB N_A2_N_c_659_n 0.0153869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A2_N_c_660_n 0.0153689f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.465
cc_129 VPB N_A2_N_c_661_n 0.0186154f $X=-0.19 $Y=1.655 $X2=1.445 $Y2=2.465
cc_130 VPB N_A2_N_c_655_n 0.0228518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_736_n 0.0146675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_737_n 0.00786211f $X=-0.19 $Y=1.655 $X2=3.625 $Y2=2.465
cc_133 VPB N_VPWR_c_738_n 4.09336e-19 $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.51
cc_134 VPB N_VPWR_c_739_n 0.00252657f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.51
cc_135 VPB N_VPWR_c_740_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.95
cc_136 VPB N_VPWR_c_741_n 0.00176953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_742_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.51
cc_138 VPB N_VPWR_c_743_n 0.00174197f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=1.51
cc_139 VPB N_VPWR_c_744_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=3.645 $Y2=1.51
cc_140 VPB N_VPWR_c_745_n 0.0133701f $X=-0.19 $Y=1.655 $X2=1.415 $Y2=2.04
cc_141 VPB N_VPWR_c_746_n 0.0408143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_747_n 0.0536098f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=2.04
cc_143 VPB N_VPWR_c_748_n 0.00452497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_749_n 0.012266f $X=-0.19 $Y=1.655 $X2=1.235 $Y2=1.95
cc_145 VPB N_VPWR_c_750_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_751_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_752_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=1.95
cc_148 VPB N_VPWR_c_753_n 0.0158018f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=2.04
cc_149 VPB N_VPWR_c_754_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_755_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_756_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_757_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_758_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_759_n 0.0105312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_760_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_761_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_735_n 0.0545663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_132_367#_c_895_n 0.001734f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.465
cc_159 VPB N_Y_c_936_n 7.8337e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_Y_c_940_n 0.00511328f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=1.535
cc_161 VPB N_Y_c_941_n 0.0027472f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 N_B1_M1034_g N_B2_M1010_g 0.0218273f $X=1.375 $Y=0.745 $X2=0 $Y2=0
cc_163 N_B1_M1036_g N_B2_M1005_g 0.0324214f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_164 B1 N_B2_M1005_g 9.29696e-19 $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_165 N_B1_c_179_p N_B2_M1005_g 0.0132999f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_166 N_B1_c_179_p N_B2_M1021_g 0.010883f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_167 N_B1_c_179_p N_B2_M1032_g 0.010883f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_168 N_B1_M1039_g N_B2_M1030_g 0.0219813f $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_169 N_B1_c_168_n N_B2_M1030_g 0.00244046f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_170 N_B1_M1038_g N_B2_M1037_g 0.0539347f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B1_c_175_n N_B2_M1037_g 0.00451525f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_172 N_B1_c_179_p N_B2_M1037_g 0.0127214f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_173 N_B1_c_187_p B2 0.0186916f $X=1.235 $Y=1.645 $X2=0 $Y2=0
cc_174 B1 B2 0.0108145f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_175 N_B1_c_167_n B2 0.00294134f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_176 N_B1_c_168_n B2 7.8499e-19 $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_177 N_B1_c_175_n B2 0.019562f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_178 N_B1_c_179_p B2 0.108608f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_179 N_B1_c_167_n N_B2_c_290_n 0.023145f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_180 N_B1_c_168_n N_B2_c_290_n 0.0226895f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_181 N_B1_c_175_n N_B2_c_290_n 0.00105603f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_182 N_B1_c_179_p N_B2_c_290_n 0.00203474f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_183 N_B1_M1039_g N_A_804_39#_M1011_g 0.0244286f $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_184 N_B1_c_168_n N_A_804_39#_M1011_g 0.023851f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_185 N_B1_M1038_g N_A_804_39#_M1002_g 0.0465537f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_186 B1 N_A_804_39#_M1002_g 7.18195e-19 $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_187 N_B1_c_175_n N_A_804_39#_M1002_g 9.60299e-19 $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_188 N_B1_c_175_n N_A_804_39#_c_377_n 2.95973e-19 $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_189 B1 N_VPWR_M1012_d 0.00206498f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_190 B1 N_VPWR_M1038_d 0.00222062f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_191 N_B1_c_175_n N_VPWR_M1038_d 9.7337e-19 $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_192 N_B1_M1009_g N_VPWR_c_737_n 0.00739639f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_193 N_B1_c_166_n N_VPWR_c_737_n 0.00566195f $X=1.055 $Y=1.535 $X2=0 $Y2=0
cc_194 N_B1_c_167_n N_VPWR_c_737_n 0.00180516f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_195 N_B1_M1009_g N_VPWR_c_738_n 5.83024e-19 $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_196 N_B1_M1012_g N_VPWR_c_738_n 0.00937807f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_197 N_B1_M1036_g N_VPWR_c_738_n 0.0105249f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_198 N_B1_M1038_g N_VPWR_c_739_n 0.00299776f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_199 N_B1_M1036_g N_VPWR_c_747_n 0.00486043f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B1_M1038_g N_VPWR_c_747_n 0.00421658f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_201 N_B1_M1009_g N_VPWR_c_753_n 0.00585385f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B1_M1012_g N_VPWR_c_753_n 0.00486043f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B1_M1009_g N_VPWR_c_735_n 0.011612f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B1_M1012_g N_VPWR_c_735_n 0.00447879f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B1_M1036_g N_VPWR_c_735_n 0.00457504f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B1_M1038_g N_VPWR_c_735_n 0.00590756f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B1_c_179_p N_A_132_367#_M1036_s 0.00484401f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_208 N_B1_c_179_p N_A_132_367#_M1021_s 0.00334892f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_209 N_B1_c_175_n N_A_132_367#_M1037_s 0.00147394f $X=3.645 $Y=1.51 $X2=0
+ $Y2=0
cc_210 N_B1_c_179_p N_A_132_367#_M1037_s 0.00746253f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_211 N_B1_M1009_g N_A_132_367#_c_895_n 4.44313e-19 $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_B1_M1012_g N_A_132_367#_c_895_n 4.11899e-19 $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_213 N_B1_c_166_n N_A_132_367#_c_895_n 0.0154288f $X=1.055 $Y=1.535 $X2=0
+ $Y2=0
cc_214 B1 N_A_132_367#_c_895_n 0.00582246f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_215 N_B1_c_167_n N_A_132_367#_c_895_n 0.00270061f $X=1.445 $Y=1.51 $X2=0
+ $Y2=0
cc_216 N_B1_M1012_g N_A_132_367#_c_905_n 0.0131492f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_217 N_B1_M1036_g N_A_132_367#_c_905_n 0.00989433f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_218 B1 N_A_132_367#_c_905_n 0.0160831f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_219 N_B1_c_167_n N_A_132_367#_c_905_n 2.82388e-19 $X=1.445 $Y=1.51 $X2=0
+ $Y2=0
cc_220 N_B1_c_179_p N_A_132_367#_c_905_n 0.00576141f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_221 N_B1_c_179_p N_A_132_367#_c_910_n 0.0132165f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_222 N_B1_M1038_g N_A_132_367#_c_911_n 0.00333139f $X=3.625 $Y=2.465 $X2=0
+ $Y2=0
cc_223 N_B1_c_179_p N_A_132_367#_c_911_n 0.00335726f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_224 N_B1_c_179_p N_Y_M1005_d 0.00334892f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_225 N_B1_c_179_p N_Y_M1032_d 0.00334892f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_226 N_B1_M1039_g N_Y_c_936_n 9.73668e-19 $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_227 N_B1_M1038_g N_Y_c_936_n 2.90083e-19 $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_228 N_B1_c_168_n N_Y_c_936_n 0.00392953f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_229 N_B1_c_175_n N_Y_c_936_n 0.0254694f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_230 N_B1_M1039_g N_Y_c_938_n 3.02451e-19 $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_231 N_B1_M1038_g N_Y_c_941_n 2.72716e-19 $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_232 N_B1_c_175_n N_Y_c_941_n 0.00911323f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_233 N_B1_M1038_g Y 0.0182666f $X=3.625 $Y=2.465 $X2=0 $Y2=0
cc_234 B1 Y 0.017555f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_235 N_B1_c_168_n Y 3.99787e-19 $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_236 N_B1_c_179_p Y 0.0820755f $X=3.48 $Y=2.04 $X2=0 $Y2=0
cc_237 N_B1_M1017_g N_A_35_65#_c_1021_n 0.0035087f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_238 N_B1_M1017_g N_A_35_65#_c_1022_n 0.0143619f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_239 N_B1_M1019_g N_A_35_65#_c_1022_n 0.0136351f $X=0.945 $Y=0.745 $X2=0 $Y2=0
cc_240 N_B1_c_166_n N_A_35_65#_c_1022_n 0.0464306f $X=1.055 $Y=1.535 $X2=0 $Y2=0
cc_241 N_B1_c_187_p N_A_35_65#_c_1022_n 7.66803e-19 $X=1.235 $Y=1.645 $X2=0
+ $Y2=0
cc_242 N_B1_c_167_n N_A_35_65#_c_1022_n 0.00363287f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_243 N_B1_M1019_g N_A_35_65#_c_1024_n 9.14714e-19 $X=0.945 $Y=0.745 $X2=0
+ $Y2=0
cc_244 N_B1_M1034_g N_A_35_65#_c_1024_n 9.14714e-19 $X=1.375 $Y=0.745 $X2=0
+ $Y2=0
cc_245 N_B1_M1034_g N_A_35_65#_c_1025_n 0.014659f $X=1.375 $Y=0.745 $X2=0 $Y2=0
cc_246 N_B1_c_187_p N_A_35_65#_c_1025_n 0.0124055f $X=1.235 $Y=1.645 $X2=0 $Y2=0
cc_247 N_B1_c_167_n N_A_35_65#_c_1025_n 0.00318714f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_248 N_B1_M1039_g N_A_35_65#_c_1029_n 0.0137525f $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_249 N_B1_c_168_n N_A_35_65#_c_1029_n 0.00511145f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_250 N_B1_c_175_n N_A_35_65#_c_1029_n 0.027095f $X=3.645 $Y=1.51 $X2=0 $Y2=0
cc_251 N_B1_M1039_g N_A_35_65#_c_1052_n 0.00310061f $X=3.605 $Y=0.745 $X2=0
+ $Y2=0
cc_252 N_B1_M1039_g N_A_35_65#_c_1053_n 0.00402124f $X=3.605 $Y=0.745 $X2=0
+ $Y2=0
cc_253 N_B1_M1039_g N_A_35_65#_c_1031_n 0.00272651f $X=3.605 $Y=0.745 $X2=0
+ $Y2=0
cc_254 N_B1_c_187_p N_A_35_65#_c_1034_n 0.0169845f $X=1.235 $Y=1.645 $X2=0 $Y2=0
cc_255 N_B1_c_167_n N_A_35_65#_c_1034_n 0.00286684f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_256 N_B1_M1039_g N_A_35_65#_c_1057_n 0.00168845f $X=3.605 $Y=0.745 $X2=0
+ $Y2=0
cc_257 N_B1_M1017_g N_VGND_c_1138_n 0.0125815f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_258 N_B1_M1019_g N_VGND_c_1138_n 0.0101212f $X=0.945 $Y=0.745 $X2=0 $Y2=0
cc_259 N_B1_M1034_g N_VGND_c_1138_n 5.09471e-19 $X=1.375 $Y=0.745 $X2=0 $Y2=0
cc_260 N_B1_M1019_g N_VGND_c_1139_n 5.09471e-19 $X=0.945 $Y=0.745 $X2=0 $Y2=0
cc_261 N_B1_M1034_g N_VGND_c_1139_n 0.0100854f $X=1.375 $Y=0.745 $X2=0 $Y2=0
cc_262 N_B1_M1039_g N_VGND_c_1141_n 0.00539667f $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_263 N_B1_M1019_g N_VGND_c_1145_n 0.00414769f $X=0.945 $Y=0.745 $X2=0 $Y2=0
cc_264 N_B1_M1034_g N_VGND_c_1145_n 0.00414769f $X=1.375 $Y=0.745 $X2=0 $Y2=0
cc_265 N_B1_M1039_g N_VGND_c_1151_n 0.00466948f $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_266 N_B1_M1017_g N_VGND_c_1153_n 0.00414769f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_267 N_B1_M1017_g N_VGND_c_1155_n 0.00824748f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_268 N_B1_M1019_g N_VGND_c_1155_n 0.00787505f $X=0.945 $Y=0.745 $X2=0 $Y2=0
cc_269 N_B1_M1034_g N_VGND_c_1155_n 0.00787505f $X=1.375 $Y=0.745 $X2=0 $Y2=0
cc_270 N_B1_M1039_g N_VGND_c_1155_n 0.00900055f $X=3.605 $Y=0.745 $X2=0 $Y2=0
cc_271 N_B2_M1005_g N_VPWR_c_738_n 0.0010486f $X=1.905 $Y=2.465 $X2=0 $Y2=0
cc_272 N_B2_M1005_g N_VPWR_c_747_n 0.00357877f $X=1.905 $Y=2.465 $X2=0 $Y2=0
cc_273 N_B2_M1021_g N_VPWR_c_747_n 0.00357877f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_274 N_B2_M1032_g N_VPWR_c_747_n 0.00357877f $X=2.765 $Y=2.465 $X2=0 $Y2=0
cc_275 N_B2_M1037_g N_VPWR_c_747_n 0.00357877f $X=3.195 $Y=2.465 $X2=0 $Y2=0
cc_276 N_B2_M1005_g N_VPWR_c_735_n 0.00544745f $X=1.905 $Y=2.465 $X2=0 $Y2=0
cc_277 N_B2_M1021_g N_VPWR_c_735_n 0.0053512f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_278 N_B2_M1032_g N_VPWR_c_735_n 0.0053512f $X=2.765 $Y=2.465 $X2=0 $Y2=0
cc_279 N_B2_M1037_g N_VPWR_c_735_n 0.00537654f $X=3.195 $Y=2.465 $X2=0 $Y2=0
cc_280 N_B2_M1005_g N_A_132_367#_c_911_n 0.0127753f $X=1.905 $Y=2.465 $X2=0
+ $Y2=0
cc_281 N_B2_M1021_g N_A_132_367#_c_911_n 0.0103812f $X=2.335 $Y=2.465 $X2=0
+ $Y2=0
cc_282 N_B2_M1032_g N_A_132_367#_c_911_n 0.0104569f $X=2.765 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_B2_M1037_g N_A_132_367#_c_911_n 0.0104569f $X=3.195 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_B2_M1021_g Y 0.0127021f $X=2.335 $Y=2.465 $X2=0 $Y2=0
cc_285 N_B2_M1032_g Y 0.0126112f $X=2.765 $Y=2.465 $X2=0 $Y2=0
cc_286 N_B2_M1037_g Y 0.0126112f $X=3.195 $Y=2.465 $X2=0 $Y2=0
cc_287 N_B2_M1010_g N_A_35_65#_c_1025_n 0.0135857f $X=1.805 $Y=0.745 $X2=0 $Y2=0
cc_288 B2 N_A_35_65#_c_1025_n 0.025009f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_289 N_B2_M1010_g N_A_35_65#_c_1026_n 8.28776e-19 $X=1.805 $Y=0.745 $X2=0
+ $Y2=0
cc_290 N_B2_M1015_g N_A_35_65#_c_1026_n 8.28776e-19 $X=2.235 $Y=0.745 $X2=0
+ $Y2=0
cc_291 N_B2_M1015_g N_A_35_65#_c_1027_n 0.0136326f $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_292 N_B2_M1029_g N_A_35_65#_c_1027_n 0.0136351f $X=2.665 $Y=0.745 $X2=0 $Y2=0
cc_293 B2 N_A_35_65#_c_1027_n 0.0496534f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_294 N_B2_c_290_n N_A_35_65#_c_1027_n 0.00289796f $X=3.195 $Y=1.51 $X2=0 $Y2=0
cc_295 N_B2_M1029_g N_A_35_65#_c_1028_n 8.28776e-19 $X=2.665 $Y=0.745 $X2=0
+ $Y2=0
cc_296 N_B2_M1030_g N_A_35_65#_c_1028_n 8.28776e-19 $X=3.095 $Y=0.745 $X2=0
+ $Y2=0
cc_297 N_B2_M1030_g N_A_35_65#_c_1029_n 0.0137139f $X=3.095 $Y=0.745 $X2=0 $Y2=0
cc_298 B2 N_A_35_65#_c_1029_n 0.0167842f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_299 N_B2_c_290_n N_A_35_65#_c_1029_n 0.00395625f $X=3.195 $Y=1.51 $X2=0 $Y2=0
cc_300 N_B2_M1030_g N_A_35_65#_c_1053_n 5.79407e-19 $X=3.095 $Y=0.745 $X2=0
+ $Y2=0
cc_301 B2 N_A_35_65#_c_1035_n 0.0161047f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_302 N_B2_c_290_n N_A_35_65#_c_1035_n 0.00299787f $X=3.195 $Y=1.51 $X2=0 $Y2=0
cc_303 B2 N_A_35_65#_c_1036_n 0.0161047f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_304 N_B2_c_290_n N_A_35_65#_c_1036_n 0.00299787f $X=3.195 $Y=1.51 $X2=0 $Y2=0
cc_305 N_B2_M1010_g N_VGND_c_1139_n 0.0100854f $X=1.805 $Y=0.745 $X2=0 $Y2=0
cc_306 N_B2_M1015_g N_VGND_c_1139_n 5.09471e-19 $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_307 N_B2_M1010_g N_VGND_c_1140_n 5.09471e-19 $X=1.805 $Y=0.745 $X2=0 $Y2=0
cc_308 N_B2_M1015_g N_VGND_c_1140_n 0.0101212f $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_309 N_B2_M1029_g N_VGND_c_1140_n 0.0101212f $X=2.665 $Y=0.745 $X2=0 $Y2=0
cc_310 N_B2_M1030_g N_VGND_c_1140_n 5.09471e-19 $X=3.095 $Y=0.745 $X2=0 $Y2=0
cc_311 N_B2_M1029_g N_VGND_c_1141_n 5.12382e-19 $X=2.665 $Y=0.745 $X2=0 $Y2=0
cc_312 N_B2_M1030_g N_VGND_c_1141_n 0.010276f $X=3.095 $Y=0.745 $X2=0 $Y2=0
cc_313 N_B2_M1010_g N_VGND_c_1147_n 0.00414769f $X=1.805 $Y=0.745 $X2=0 $Y2=0
cc_314 N_B2_M1015_g N_VGND_c_1147_n 0.00414769f $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_315 N_B2_M1029_g N_VGND_c_1149_n 0.00414769f $X=2.665 $Y=0.745 $X2=0 $Y2=0
cc_316 N_B2_M1030_g N_VGND_c_1149_n 0.00414769f $X=3.095 $Y=0.745 $X2=0 $Y2=0
cc_317 N_B2_M1010_g N_VGND_c_1155_n 0.00787505f $X=1.805 $Y=0.745 $X2=0 $Y2=0
cc_318 N_B2_M1015_g N_VGND_c_1155_n 0.00787505f $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_319 N_B2_M1029_g N_VGND_c_1155_n 0.00787505f $X=2.665 $Y=0.745 $X2=0 $Y2=0
cc_320 N_B2_M1030_g N_VGND_c_1155_n 0.00787505f $X=3.095 $Y=0.745 $X2=0 $Y2=0
cc_321 N_A_804_39#_M1025_g N_A1_N_M1000_g 0.00631592f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_322 N_A_804_39#_c_383_n N_A1_N_M1000_g 0.014624f $X=6.28 $Y=1.855 $X2=0 $Y2=0
cc_323 N_A_804_39#_c_385_n N_A1_N_M1006_g 0.0134041f $X=7.14 $Y=1.855 $X2=0
+ $Y2=0
cc_324 N_A_804_39#_c_385_n N_A1_N_M1022_g 0.0134041f $X=7.14 $Y=1.855 $X2=0
+ $Y2=0
cc_325 N_A_804_39#_c_386_n N_A1_N_M1026_g 0.0147693f $X=8.34 $Y=1.855 $X2=0
+ $Y2=0
cc_326 N_A_804_39#_c_386_n N_A1_N_c_562_n 0.0428647f $X=8.34 $Y=1.855 $X2=0
+ $Y2=0
cc_327 N_A_804_39#_c_391_n N_A1_N_c_562_n 0.0153308f $X=7.235 $Y=1.855 $X2=0
+ $Y2=0
cc_328 N_A_804_39#_c_372_n N_A1_N_c_563_n 4.88939e-19 $X=5.555 $Y=1.51 $X2=0
+ $Y2=0
cc_329 N_A_804_39#_c_373_n N_A1_N_c_563_n 0.00315766f $X=5.64 $Y=1.765 $X2=0
+ $Y2=0
cc_330 N_A_804_39#_c_385_n N_A1_N_c_563_n 0.00279051f $X=7.14 $Y=1.855 $X2=0
+ $Y2=0
cc_331 N_A_804_39#_c_386_n N_A1_N_c_563_n 0.0112154f $X=8.34 $Y=1.855 $X2=0
+ $Y2=0
cc_332 N_A_804_39#_c_390_n N_A1_N_c_563_n 0.00256759f $X=6.375 $Y=1.855 $X2=0
+ $Y2=0
cc_333 N_A_804_39#_c_391_n N_A1_N_c_563_n 0.0028903f $X=7.235 $Y=1.855 $X2=0
+ $Y2=0
cc_334 N_A_804_39#_c_377_n N_A1_N_c_563_n 0.00972845f $X=5.565 $Y=1.51 $X2=0
+ $Y2=0
cc_335 N_A_804_39#_M1031_g N_A1_N_c_564_n 0.00435239f $X=5.565 $Y=0.745 $X2=0
+ $Y2=0
cc_336 N_A_804_39#_c_372_n N_A1_N_c_564_n 0.0151985f $X=5.555 $Y=1.51 $X2=0
+ $Y2=0
cc_337 N_A_804_39#_c_383_n N_A1_N_c_564_n 0.0287983f $X=6.28 $Y=1.855 $X2=0
+ $Y2=0
cc_338 N_A_804_39#_c_390_n N_A1_N_c_564_n 0.0161566f $X=6.375 $Y=1.855 $X2=0
+ $Y2=0
cc_339 N_A_804_39#_c_377_n N_A1_N_c_564_n 0.00297316f $X=5.565 $Y=1.51 $X2=0
+ $Y2=0
cc_340 N_A_804_39#_c_385_n N_A1_N_c_565_n 0.0473335f $X=7.14 $Y=1.855 $X2=0
+ $Y2=0
cc_341 N_A_804_39#_c_386_n N_A2_N_c_658_n 0.0190006f $X=8.34 $Y=1.855 $X2=-0.19
+ $Y2=-0.245
cc_342 N_A_804_39#_c_422_p N_A2_N_M1001_g 0.00499458f $X=8.45 $Y=0.77 $X2=0
+ $Y2=0
cc_343 N_A_804_39#_c_387_n N_A2_N_c_659_n 0.0134041f $X=9.21 $Y=1.855 $X2=0
+ $Y2=0
cc_344 N_A_804_39#_c_424_p N_A2_N_M1016_g 0.0100683f $X=9.145 $Y=0.907 $X2=0
+ $Y2=0
cc_345 N_A_804_39#_c_376_n N_A2_N_M1016_g 0.00146517f $X=9.31 $Y=0.7 $X2=0 $Y2=0
cc_346 N_A_804_39#_c_387_n N_A2_N_c_660_n 0.0134041f $X=9.21 $Y=1.855 $X2=0
+ $Y2=0
cc_347 N_A_804_39#_c_424_p N_A2_N_M1018_g 0.010826f $X=9.145 $Y=0.907 $X2=0
+ $Y2=0
cc_348 N_A_804_39#_c_376_n N_A2_N_M1018_g 0.0102056f $X=9.31 $Y=0.7 $X2=0 $Y2=0
cc_349 N_A_804_39#_c_388_n N_A2_N_c_661_n 0.0151009f $X=9.815 $Y=1.855 $X2=0
+ $Y2=0
cc_350 N_A_804_39#_c_374_n N_A2_N_M1020_g 0.0121838f $X=9.815 $Y=1.165 $X2=0
+ $Y2=0
cc_351 N_A_804_39#_c_375_n N_A2_N_M1020_g 0.00292251f $X=9.905 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A_804_39#_c_376_n N_A2_N_M1020_g 0.0133801f $X=9.31 $Y=0.7 $X2=0 $Y2=0
cc_353 N_A_804_39#_c_424_p N_A2_N_c_654_n 0.0047792f $X=9.145 $Y=0.907 $X2=0
+ $Y2=0
cc_354 N_A_804_39#_c_388_n N_A2_N_c_654_n 0.0170004f $X=9.815 $Y=1.855 $X2=0
+ $Y2=0
cc_355 N_A_804_39#_c_374_n N_A2_N_c_654_n 0.0110246f $X=9.815 $Y=1.165 $X2=0
+ $Y2=0
cc_356 N_A_804_39#_c_375_n N_A2_N_c_654_n 0.0129078f $X=9.905 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_A_804_39#_c_376_n N_A2_N_c_654_n 0.0261484f $X=9.31 $Y=0.7 $X2=0 $Y2=0
cc_358 N_A_804_39#_c_393_n N_A2_N_c_654_n 0.0145234f $X=9.3 $Y=1.855 $X2=0 $Y2=0
cc_359 N_A_804_39#_c_387_n N_A2_N_c_655_n 0.00275477f $X=9.21 $Y=1.855 $X2=0
+ $Y2=0
cc_360 N_A_804_39#_c_424_p N_A2_N_c_655_n 4.65218e-19 $X=9.145 $Y=0.907 $X2=0
+ $Y2=0
cc_361 N_A_804_39#_c_388_n N_A2_N_c_655_n 0.00129855f $X=9.815 $Y=1.855 $X2=0
+ $Y2=0
cc_362 N_A_804_39#_c_374_n N_A2_N_c_655_n 8.63852e-19 $X=9.815 $Y=1.165 $X2=0
+ $Y2=0
cc_363 N_A_804_39#_c_375_n N_A2_N_c_655_n 0.0110648f $X=9.905 $Y=1.765 $X2=0
+ $Y2=0
cc_364 N_A_804_39#_c_422_p N_A2_N_c_655_n 4.95895e-19 $X=8.45 $Y=0.77 $X2=0
+ $Y2=0
cc_365 N_A_804_39#_c_392_n N_A2_N_c_655_n 0.00286534f $X=8.435 $Y=1.855 $X2=0
+ $Y2=0
cc_366 N_A_804_39#_c_376_n N_A2_N_c_655_n 0.00268527f $X=9.31 $Y=0.7 $X2=0 $Y2=0
cc_367 N_A_804_39#_c_393_n N_A2_N_c_655_n 0.00286534f $X=9.3 $Y=1.855 $X2=0
+ $Y2=0
cc_368 N_A_804_39#_c_386_n N_A2_N_c_656_n 0.00415816f $X=8.34 $Y=1.855 $X2=0
+ $Y2=0
cc_369 N_A_804_39#_c_387_n N_A2_N_c_656_n 0.049858f $X=9.21 $Y=1.855 $X2=0 $Y2=0
cc_370 N_A_804_39#_c_424_p N_A2_N_c_656_n 0.0274448f $X=9.145 $Y=0.907 $X2=0
+ $Y2=0
cc_371 N_A_804_39#_c_422_p N_A2_N_c_656_n 0.0206472f $X=8.45 $Y=0.77 $X2=0 $Y2=0
cc_372 N_A_804_39#_c_392_n N_A2_N_c_656_n 0.0163065f $X=8.435 $Y=1.855 $X2=0
+ $Y2=0
cc_373 N_A_804_39#_c_376_n N_A2_N_c_657_n 0.00709151f $X=9.31 $Y=0.7 $X2=0 $Y2=0
cc_374 N_A_804_39#_c_383_n N_VPWR_M1025_s 0.00420909f $X=6.28 $Y=1.855 $X2=0
+ $Y2=0
cc_375 N_A_804_39#_c_384_n N_VPWR_M1025_s 0.0039124f $X=5.725 $Y=1.855 $X2=0
+ $Y2=0
cc_376 N_A_804_39#_c_385_n N_VPWR_M1006_d 0.00181066f $X=7.14 $Y=1.855 $X2=0
+ $Y2=0
cc_377 N_A_804_39#_c_386_n N_VPWR_M1026_d 0.00708787f $X=8.34 $Y=1.855 $X2=0
+ $Y2=0
cc_378 N_A_804_39#_c_387_n N_VPWR_M1014_s 0.00181066f $X=9.21 $Y=1.855 $X2=0
+ $Y2=0
cc_379 N_A_804_39#_c_388_n N_VPWR_M1033_s 0.00272766f $X=9.815 $Y=1.855 $X2=0
+ $Y2=0
cc_380 N_A_804_39#_M1002_g N_VPWR_c_739_n 0.00695533f $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_381 N_A_804_39#_M1008_g N_VPWR_c_739_n 5.25742e-19 $X=4.525 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_A_804_39#_M1002_g N_VPWR_c_740_n 7.52785e-19 $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_383 N_A_804_39#_M1008_g N_VPWR_c_740_n 0.0140093f $X=4.525 $Y=2.465 $X2=0
+ $Y2=0
cc_384 N_A_804_39#_M1013_g N_VPWR_c_740_n 0.0140168f $X=4.955 $Y=2.465 $X2=0
+ $Y2=0
cc_385 N_A_804_39#_M1025_g N_VPWR_c_740_n 7.21513e-19 $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_A_804_39#_M1013_g N_VPWR_c_741_n 7.31032e-19 $X=4.955 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_A_804_39#_M1025_g N_VPWR_c_741_n 0.0152068f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_A_804_39#_c_372_n N_VPWR_c_741_n 0.00269032f $X=5.555 $Y=1.51 $X2=0
+ $Y2=0
cc_389 N_A_804_39#_c_383_n N_VPWR_c_741_n 0.0253884f $X=6.28 $Y=1.855 $X2=0
+ $Y2=0
cc_390 N_A_804_39#_c_384_n N_VPWR_c_741_n 0.0143958f $X=5.725 $Y=1.855 $X2=0
+ $Y2=0
cc_391 N_A_804_39#_c_377_n N_VPWR_c_741_n 0.00252906f $X=5.565 $Y=1.51 $X2=0
+ $Y2=0
cc_392 N_A_804_39#_c_385_n N_VPWR_c_742_n 0.0164152f $X=7.14 $Y=1.855 $X2=0
+ $Y2=0
cc_393 N_A_804_39#_c_386_n N_VPWR_c_743_n 0.0430217f $X=8.34 $Y=1.855 $X2=0
+ $Y2=0
cc_394 N_A_804_39#_c_387_n N_VPWR_c_744_n 0.0164152f $X=9.21 $Y=1.855 $X2=0
+ $Y2=0
cc_395 N_A_804_39#_c_388_n N_VPWR_c_746_n 0.0226958f $X=9.815 $Y=1.855 $X2=0
+ $Y2=0
cc_396 N_A_804_39#_M1002_g N_VPWR_c_749_n 0.00361126f $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_A_804_39#_M1008_g N_VPWR_c_749_n 0.00486043f $X=4.525 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_A_804_39#_c_478_p N_VPWR_c_751_n 0.0124525f $X=6.375 $Y=1.98 $X2=0
+ $Y2=0
cc_399 N_A_804_39#_M1013_g N_VPWR_c_754_n 0.00486043f $X=4.955 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A_804_39#_M1025_g N_VPWR_c_754_n 0.00486043f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_804_39#_c_481_p N_VPWR_c_755_n 0.0124525f $X=7.235 $Y=1.98 $X2=0
+ $Y2=0
cc_402 N_A_804_39#_c_482_p N_VPWR_c_756_n 0.0124525f $X=8.435 $Y=1.98 $X2=0
+ $Y2=0
cc_403 N_A_804_39#_c_483_p N_VPWR_c_757_n 0.0120977f $X=9.295 $Y=1.98 $X2=0
+ $Y2=0
cc_404 N_A_804_39#_M1000_s N_VPWR_c_735_n 0.00536646f $X=6.235 $Y=1.835 $X2=0
+ $Y2=0
cc_405 N_A_804_39#_M1022_s N_VPWR_c_735_n 0.00536646f $X=7.095 $Y=1.835 $X2=0
+ $Y2=0
cc_406 N_A_804_39#_M1007_d N_VPWR_c_735_n 0.00536646f $X=8.295 $Y=1.835 $X2=0
+ $Y2=0
cc_407 N_A_804_39#_M1028_d N_VPWR_c_735_n 0.00571434f $X=9.155 $Y=1.835 $X2=0
+ $Y2=0
cc_408 N_A_804_39#_M1002_g N_VPWR_c_735_n 0.00424777f $X=4.095 $Y=2.465 $X2=0
+ $Y2=0
cc_409 N_A_804_39#_M1008_g N_VPWR_c_735_n 0.00824727f $X=4.525 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_A_804_39#_M1013_g N_VPWR_c_735_n 0.00824727f $X=4.955 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A_804_39#_M1025_g N_VPWR_c_735_n 0.00824727f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A_804_39#_c_478_p N_VPWR_c_735_n 0.00730901f $X=6.375 $Y=1.98 $X2=0
+ $Y2=0
cc_413 N_A_804_39#_c_481_p N_VPWR_c_735_n 0.00730901f $X=7.235 $Y=1.98 $X2=0
+ $Y2=0
cc_414 N_A_804_39#_c_482_p N_VPWR_c_735_n 0.00730901f $X=8.435 $Y=1.98 $X2=0
+ $Y2=0
cc_415 N_A_804_39#_c_483_p N_VPWR_c_735_n 0.00691495f $X=9.295 $Y=1.98 $X2=0
+ $Y2=0
cc_416 N_A_804_39#_M1011_g N_Y_c_936_n 0.00230877f $X=4.095 $Y=0.745 $X2=0 $Y2=0
cc_417 N_A_804_39#_M1002_g N_Y_c_936_n 0.00240661f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_418 N_A_804_39#_M1008_g N_Y_c_936_n 3.06683e-19 $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_419 N_A_804_39#_M1023_g N_Y_c_936_n 3.02009e-19 $X=4.545 $Y=0.745 $X2=0 $Y2=0
cc_420 N_A_804_39#_c_372_n N_Y_c_936_n 0.0122207f $X=5.555 $Y=1.51 $X2=0 $Y2=0
cc_421 N_A_804_39#_c_377_n N_Y_c_936_n 0.0146406f $X=5.565 $Y=1.51 $X2=0 $Y2=0
cc_422 N_A_804_39#_M1002_g N_Y_c_964_n 0.00720543f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_423 N_A_804_39#_M1011_g N_Y_c_965_n 0.00486574f $X=4.095 $Y=0.745 $X2=0 $Y2=0
cc_424 N_A_804_39#_M1023_g N_Y_c_965_n 0.00684536f $X=4.545 $Y=0.745 $X2=0 $Y2=0
cc_425 N_A_804_39#_M1027_g N_Y_c_965_n 6.31572e-19 $X=5.055 $Y=0.745 $X2=0 $Y2=0
cc_426 N_A_804_39#_M1008_g N_Y_c_940_n 0.0129702f $X=4.525 $Y=2.465 $X2=0 $Y2=0
cc_427 N_A_804_39#_M1013_g N_Y_c_940_n 0.0128776f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_428 N_A_804_39#_M1025_g N_Y_c_940_n 6.33061e-19 $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_429 N_A_804_39#_c_372_n N_Y_c_940_n 0.0593934f $X=5.555 $Y=1.51 $X2=0 $Y2=0
cc_430 N_A_804_39#_c_384_n N_Y_c_940_n 0.00715935f $X=5.725 $Y=1.855 $X2=0 $Y2=0
cc_431 N_A_804_39#_c_377_n N_Y_c_940_n 0.00551486f $X=5.565 $Y=1.51 $X2=0 $Y2=0
cc_432 N_A_804_39#_M1023_g N_Y_c_937_n 0.00965873f $X=4.545 $Y=0.745 $X2=0 $Y2=0
cc_433 N_A_804_39#_M1027_g N_Y_c_937_n 0.0132524f $X=5.055 $Y=0.745 $X2=0 $Y2=0
cc_434 N_A_804_39#_M1031_g N_Y_c_937_n 0.00847302f $X=5.565 $Y=0.745 $X2=0 $Y2=0
cc_435 N_A_804_39#_c_372_n N_Y_c_937_n 0.0714016f $X=5.555 $Y=1.51 $X2=0 $Y2=0
cc_436 N_A_804_39#_c_377_n N_Y_c_937_n 0.0101788f $X=5.565 $Y=1.51 $X2=0 $Y2=0
cc_437 N_A_804_39#_M1031_g N_Y_c_979_n 0.00633842f $X=5.565 $Y=0.745 $X2=0 $Y2=0
cc_438 N_A_804_39#_M1011_g N_Y_c_938_n 0.00861061f $X=4.095 $Y=0.745 $X2=0 $Y2=0
cc_439 N_A_804_39#_M1023_g N_Y_c_938_n 0.00172515f $X=4.545 $Y=0.745 $X2=0 $Y2=0
cc_440 N_A_804_39#_c_372_n N_Y_c_938_n 0.0114223f $X=5.555 $Y=1.51 $X2=0 $Y2=0
cc_441 N_A_804_39#_c_377_n N_Y_c_938_n 0.00361308f $X=5.565 $Y=1.51 $X2=0 $Y2=0
cc_442 N_A_804_39#_M1002_g N_Y_c_941_n 0.00400407f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_443 N_A_804_39#_c_372_n N_Y_c_941_n 0.0046385f $X=5.555 $Y=1.51 $X2=0 $Y2=0
cc_444 N_A_804_39#_c_377_n N_Y_c_941_n 0.00304159f $X=5.565 $Y=1.51 $X2=0 $Y2=0
cc_445 N_A_804_39#_M1002_g Y 0.0123228f $X=4.095 $Y=2.465 $X2=0 $Y2=0
cc_446 N_A_804_39#_M1011_g N_A_35_65#_c_1029_n 6.72584e-19 $X=4.095 $Y=0.745
+ $X2=0 $Y2=0
cc_447 N_A_804_39#_M1011_g N_A_35_65#_c_1053_n 0.00133027f $X=4.095 $Y=0.745
+ $X2=0 $Y2=0
cc_448 N_A_804_39#_M1011_g N_A_35_65#_c_1030_n 0.0119025f $X=4.095 $Y=0.745
+ $X2=0 $Y2=0
cc_449 N_A_804_39#_M1023_g N_A_35_65#_c_1030_n 0.0118301f $X=4.545 $Y=0.745
+ $X2=0 $Y2=0
cc_450 N_A_804_39#_M1027_g N_A_35_65#_c_1080_n 0.00675522f $X=5.055 $Y=0.745
+ $X2=0 $Y2=0
cc_451 N_A_804_39#_M1031_g N_A_35_65#_c_1080_n 5.84315e-19 $X=5.565 $Y=0.745
+ $X2=0 $Y2=0
cc_452 N_A_804_39#_M1027_g N_A_35_65#_c_1032_n 0.00875863f $X=5.055 $Y=0.745
+ $X2=0 $Y2=0
cc_453 N_A_804_39#_M1031_g N_A_35_65#_c_1032_n 0.0128765f $X=5.565 $Y=0.745
+ $X2=0 $Y2=0
cc_454 N_A_804_39#_c_372_n N_A_35_65#_c_1033_n 0.00164064f $X=5.555 $Y=1.51
+ $X2=0 $Y2=0
cc_455 N_A_804_39#_M1027_g N_A_35_65#_c_1037_n 0.00141323f $X=5.055 $Y=0.745
+ $X2=0 $Y2=0
cc_456 N_A_804_39#_M1011_g N_VGND_c_1151_n 0.0030414f $X=4.095 $Y=0.745 $X2=0
+ $Y2=0
cc_457 N_A_804_39#_M1023_g N_VGND_c_1151_n 0.0030414f $X=4.545 $Y=0.745 $X2=0
+ $Y2=0
cc_458 N_A_804_39#_M1027_g N_VGND_c_1151_n 0.00304113f $X=5.055 $Y=0.745 $X2=0
+ $Y2=0
cc_459 N_A_804_39#_M1031_g N_VGND_c_1151_n 0.0030414f $X=5.565 $Y=0.745 $X2=0
+ $Y2=0
cc_460 N_A_804_39#_M1011_g N_VGND_c_1155_n 0.00439456f $X=4.095 $Y=0.745 $X2=0
+ $Y2=0
cc_461 N_A_804_39#_M1023_g N_VGND_c_1155_n 0.00444263f $X=4.545 $Y=0.745 $X2=0
+ $Y2=0
cc_462 N_A_804_39#_M1027_g N_VGND_c_1155_n 0.0044974f $X=5.055 $Y=0.745 $X2=0
+ $Y2=0
cc_463 N_A_804_39#_M1031_g N_VGND_c_1155_n 0.0049228f $X=5.565 $Y=0.745 $X2=0
+ $Y2=0
cc_464 N_A_804_39#_c_424_p N_VGND_c_1155_n 0.00128659f $X=9.145 $Y=0.907 $X2=0
+ $Y2=0
cc_465 N_A_804_39#_c_424_p N_A_1235_65#_M1016_d 0.00338621f $X=9.145 $Y=0.907
+ $X2=0 $Y2=0
cc_466 N_A_804_39#_c_374_n N_A_1235_65#_M1020_d 0.00392559f $X=9.815 $Y=1.165
+ $X2=0 $Y2=0
cc_467 N_A_804_39#_M1031_g N_A_1235_65#_c_1274_n 2.35901e-19 $X=5.565 $Y=0.745
+ $X2=0 $Y2=0
cc_468 N_A_804_39#_c_386_n N_A_1235_65#_c_1276_n 0.00701811f $X=8.34 $Y=1.855
+ $X2=0 $Y2=0
cc_469 N_A_804_39#_M1001_s N_A_1235_65#_c_1277_n 0.00176461f $X=8.31 $Y=0.325
+ $X2=0 $Y2=0
cc_470 N_A_804_39#_c_424_p N_A_1235_65#_c_1277_n 0.00459988f $X=9.145 $Y=0.907
+ $X2=0 $Y2=0
cc_471 N_A_804_39#_c_422_p N_A_1235_65#_c_1277_n 0.0137588f $X=8.45 $Y=0.77
+ $X2=0 $Y2=0
cc_472 N_A_804_39#_M1018_s N_A_1235_65#_c_1279_n 0.00176461f $X=9.17 $Y=0.325
+ $X2=0 $Y2=0
cc_473 N_A_804_39#_c_424_p N_A_1235_65#_c_1279_n 0.00384121f $X=9.145 $Y=0.907
+ $X2=0 $Y2=0
cc_474 N_A_804_39#_c_374_n N_A_1235_65#_c_1279_n 0.0028241f $X=9.815 $Y=1.165
+ $X2=0 $Y2=0
cc_475 N_A_804_39#_c_376_n N_A_1235_65#_c_1279_n 0.0159589f $X=9.31 $Y=0.7 $X2=0
+ $Y2=0
cc_476 N_A_804_39#_c_374_n N_A_1235_65#_c_1280_n 0.0281102f $X=9.815 $Y=1.165
+ $X2=0 $Y2=0
cc_477 N_A_804_39#_c_424_p N_A_1235_65#_c_1282_n 0.0120271f $X=9.145 $Y=0.907
+ $X2=0 $Y2=0
cc_478 N_A1_N_M1035_g N_A2_N_M1001_g 0.0198152f $X=7.805 $Y=0.745 $X2=0 $Y2=0
cc_479 N_A1_N_M1026_g N_A2_N_c_655_n 0.00799346f $X=7.45 $Y=2.465 $X2=0 $Y2=0
cc_480 N_A1_N_c_562_n N_A2_N_c_655_n 7.47556e-19 $X=7.77 $Y=1.51 $X2=0 $Y2=0
cc_481 N_A1_N_c_563_n N_A2_N_c_655_n 0.0230747f $X=7.805 $Y=1.51 $X2=0 $Y2=0
cc_482 N_A1_N_M1035_g N_A2_N_c_656_n 5.34464e-19 $X=7.805 $Y=0.745 $X2=0 $Y2=0
cc_483 N_A1_N_c_562_n N_A2_N_c_656_n 0.00792948f $X=7.77 $Y=1.51 $X2=0 $Y2=0
cc_484 N_A1_N_c_563_n N_A2_N_c_656_n 6.42529e-19 $X=7.805 $Y=1.51 $X2=0 $Y2=0
cc_485 N_A1_N_M1000_g N_VPWR_c_741_n 0.0149244f $X=6.16 $Y=2.465 $X2=0 $Y2=0
cc_486 N_A1_N_M1006_g N_VPWR_c_741_n 7.31032e-19 $X=6.59 $Y=2.465 $X2=0 $Y2=0
cc_487 N_A1_N_M1000_g N_VPWR_c_742_n 7.18684e-19 $X=6.16 $Y=2.465 $X2=0 $Y2=0
cc_488 N_A1_N_M1006_g N_VPWR_c_742_n 0.0139258f $X=6.59 $Y=2.465 $X2=0 $Y2=0
cc_489 N_A1_N_M1022_g N_VPWR_c_742_n 0.0139258f $X=7.02 $Y=2.465 $X2=0 $Y2=0
cc_490 N_A1_N_M1026_g N_VPWR_c_742_n 7.18684e-19 $X=7.45 $Y=2.465 $X2=0 $Y2=0
cc_491 N_A1_N_M1022_g N_VPWR_c_743_n 7.30895e-19 $X=7.02 $Y=2.465 $X2=0 $Y2=0
cc_492 N_A1_N_M1026_g N_VPWR_c_743_n 0.0149151f $X=7.45 $Y=2.465 $X2=0 $Y2=0
cc_493 N_A1_N_M1000_g N_VPWR_c_751_n 0.00486043f $X=6.16 $Y=2.465 $X2=0 $Y2=0
cc_494 N_A1_N_M1006_g N_VPWR_c_751_n 0.00486043f $X=6.59 $Y=2.465 $X2=0 $Y2=0
cc_495 N_A1_N_M1022_g N_VPWR_c_755_n 0.00486043f $X=7.02 $Y=2.465 $X2=0 $Y2=0
cc_496 N_A1_N_M1026_g N_VPWR_c_755_n 0.00486043f $X=7.45 $Y=2.465 $X2=0 $Y2=0
cc_497 N_A1_N_M1000_g N_VPWR_c_735_n 0.00824727f $X=6.16 $Y=2.465 $X2=0 $Y2=0
cc_498 N_A1_N_M1006_g N_VPWR_c_735_n 0.00824727f $X=6.59 $Y=2.465 $X2=0 $Y2=0
cc_499 N_A1_N_M1022_g N_VPWR_c_735_n 0.00824727f $X=7.02 $Y=2.465 $X2=0 $Y2=0
cc_500 N_A1_N_M1026_g N_VPWR_c_735_n 0.00824727f $X=7.45 $Y=2.465 $X2=0 $Y2=0
cc_501 N_A1_N_c_564_n N_Y_c_937_n 0.00162095f $X=6.373 $Y=1.402 $X2=0 $Y2=0
cc_502 N_A1_N_M1003_g N_A_35_65#_c_1032_n 9.35491e-19 $X=6.515 $Y=0.745 $X2=0
+ $Y2=0
cc_503 N_A1_N_c_564_n N_A_35_65#_c_1033_n 0.00348845f $X=6.373 $Y=1.402 $X2=0
+ $Y2=0
cc_504 N_A1_N_M1003_g N_VGND_c_1142_n 0.010097f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_505 N_A1_N_M1004_g N_VGND_c_1142_n 0.00878393f $X=6.945 $Y=0.745 $X2=0 $Y2=0
cc_506 N_A1_N_M1024_g N_VGND_c_1142_n 4.51475e-19 $X=7.375 $Y=0.745 $X2=0 $Y2=0
cc_507 N_A1_N_M1004_g N_VGND_c_1143_n 0.00414769f $X=6.945 $Y=0.745 $X2=0 $Y2=0
cc_508 N_A1_N_M1024_g N_VGND_c_1143_n 0.00414769f $X=7.375 $Y=0.745 $X2=0 $Y2=0
cc_509 N_A1_N_M1004_g N_VGND_c_1144_n 4.99852e-19 $X=6.945 $Y=0.745 $X2=0 $Y2=0
cc_510 N_A1_N_M1024_g N_VGND_c_1144_n 0.0101212f $X=7.375 $Y=0.745 $X2=0 $Y2=0
cc_511 N_A1_N_M1035_g N_VGND_c_1144_n 0.0102472f $X=7.805 $Y=0.745 $X2=0 $Y2=0
cc_512 N_A1_N_M1003_g N_VGND_c_1151_n 0.00414769f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_513 N_A1_N_M1035_g N_VGND_c_1154_n 0.00414769f $X=7.805 $Y=0.745 $X2=0 $Y2=0
cc_514 N_A1_N_M1003_g N_VGND_c_1155_n 0.00837493f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_515 N_A1_N_M1004_g N_VGND_c_1155_n 0.00787505f $X=6.945 $Y=0.745 $X2=0 $Y2=0
cc_516 N_A1_N_M1024_g N_VGND_c_1155_n 0.00787505f $X=7.375 $Y=0.745 $X2=0 $Y2=0
cc_517 N_A1_N_M1035_g N_VGND_c_1155_n 0.0078848f $X=7.805 $Y=0.745 $X2=0 $Y2=0
cc_518 N_A1_N_c_563_n N_A_1235_65#_c_1273_n 0.00145819f $X=7.805 $Y=1.51 $X2=0
+ $Y2=0
cc_519 N_A1_N_c_564_n N_A_1235_65#_c_1273_n 0.022285f $X=6.373 $Y=1.402 $X2=0
+ $Y2=0
cc_520 N_A1_N_M1003_g N_A_1235_65#_c_1274_n 0.0022867f $X=6.515 $Y=0.745 $X2=0
+ $Y2=0
cc_521 N_A1_N_M1003_g N_A_1235_65#_c_1299_n 0.0122209f $X=6.515 $Y=0.745 $X2=0
+ $Y2=0
cc_522 N_A1_N_M1004_g N_A_1235_65#_c_1299_n 0.013248f $X=6.945 $Y=0.745 $X2=0
+ $Y2=0
cc_523 N_A1_N_c_562_n N_A_1235_65#_c_1299_n 0.0149439f $X=7.77 $Y=1.51 $X2=0
+ $Y2=0
cc_524 N_A1_N_c_563_n N_A_1235_65#_c_1299_n 0.00236086f $X=7.805 $Y=1.51 $X2=0
+ $Y2=0
cc_525 N_A1_N_c_565_n N_A_1235_65#_c_1299_n 0.0109224f $X=6.565 $Y=1.402 $X2=0
+ $Y2=0
cc_526 N_A1_N_M1004_g N_A_1235_65#_c_1275_n 8.28776e-19 $X=6.945 $Y=0.745 $X2=0
+ $Y2=0
cc_527 N_A1_N_M1024_g N_A_1235_65#_c_1275_n 8.28776e-19 $X=7.375 $Y=0.745 $X2=0
+ $Y2=0
cc_528 N_A1_N_M1024_g N_A_1235_65#_c_1276_n 0.0126391f $X=7.375 $Y=0.745 $X2=0
+ $Y2=0
cc_529 N_A1_N_M1035_g N_A_1235_65#_c_1276_n 0.0130183f $X=7.805 $Y=0.745 $X2=0
+ $Y2=0
cc_530 N_A1_N_c_562_n N_A_1235_65#_c_1276_n 0.0455144f $X=7.77 $Y=1.51 $X2=0
+ $Y2=0
cc_531 N_A1_N_c_563_n N_A_1235_65#_c_1276_n 0.00380394f $X=7.805 $Y=1.51 $X2=0
+ $Y2=0
cc_532 N_A1_N_M1035_g N_A_1235_65#_c_1278_n 4.90985e-19 $X=7.805 $Y=0.745 $X2=0
+ $Y2=0
cc_533 N_A1_N_M1004_g N_A_1235_65#_c_1281_n 0.00154451f $X=6.945 $Y=0.745 $X2=0
+ $Y2=0
cc_534 N_A1_N_c_562_n N_A_1235_65#_c_1281_n 0.015271f $X=7.77 $Y=1.51 $X2=0
+ $Y2=0
cc_535 N_A1_N_c_563_n N_A_1235_65#_c_1281_n 0.00287441f $X=7.805 $Y=1.51 $X2=0
+ $Y2=0
cc_536 N_A1_N_c_565_n N_A_1235_65#_c_1281_n 0.00122552f $X=6.565 $Y=1.402 $X2=0
+ $Y2=0
cc_537 N_A2_N_c_658_n N_VPWR_c_743_n 0.0149151f $X=8.22 $Y=1.725 $X2=0 $Y2=0
cc_538 N_A2_N_c_659_n N_VPWR_c_743_n 7.30895e-19 $X=8.65 $Y=1.725 $X2=0 $Y2=0
cc_539 N_A2_N_c_658_n N_VPWR_c_744_n 7.18684e-19 $X=8.22 $Y=1.725 $X2=0 $Y2=0
cc_540 N_A2_N_c_659_n N_VPWR_c_744_n 0.0139258f $X=8.65 $Y=1.725 $X2=0 $Y2=0
cc_541 N_A2_N_c_660_n N_VPWR_c_744_n 0.0141441f $X=9.08 $Y=1.725 $X2=0 $Y2=0
cc_542 N_A2_N_c_661_n N_VPWR_c_744_n 7.33419e-19 $X=9.51 $Y=1.725 $X2=0 $Y2=0
cc_543 N_A2_N_c_660_n N_VPWR_c_746_n 7.21513e-19 $X=9.08 $Y=1.725 $X2=0 $Y2=0
cc_544 N_A2_N_c_661_n N_VPWR_c_746_n 0.0150803f $X=9.51 $Y=1.725 $X2=0 $Y2=0
cc_545 N_A2_N_c_658_n N_VPWR_c_756_n 0.00486043f $X=8.22 $Y=1.725 $X2=0 $Y2=0
cc_546 N_A2_N_c_659_n N_VPWR_c_756_n 0.00486043f $X=8.65 $Y=1.725 $X2=0 $Y2=0
cc_547 N_A2_N_c_660_n N_VPWR_c_757_n 0.00486043f $X=9.08 $Y=1.725 $X2=0 $Y2=0
cc_548 N_A2_N_c_661_n N_VPWR_c_757_n 0.00486043f $X=9.51 $Y=1.725 $X2=0 $Y2=0
cc_549 N_A2_N_c_658_n N_VPWR_c_735_n 0.00824727f $X=8.22 $Y=1.725 $X2=0 $Y2=0
cc_550 N_A2_N_c_659_n N_VPWR_c_735_n 0.00824727f $X=8.65 $Y=1.725 $X2=0 $Y2=0
cc_551 N_A2_N_c_660_n N_VPWR_c_735_n 0.00824727f $X=9.08 $Y=1.725 $X2=0 $Y2=0
cc_552 N_A2_N_c_661_n N_VPWR_c_735_n 0.00824727f $X=9.51 $Y=1.725 $X2=0 $Y2=0
cc_553 N_A2_N_M1001_g N_VGND_c_1144_n 5.59621e-19 $X=8.235 $Y=0.745 $X2=0 $Y2=0
cc_554 N_A2_N_M1001_g N_VGND_c_1154_n 0.0030414f $X=8.235 $Y=0.745 $X2=0 $Y2=0
cc_555 N_A2_N_M1016_g N_VGND_c_1154_n 0.0030414f $X=8.665 $Y=0.745 $X2=0 $Y2=0
cc_556 N_A2_N_M1018_g N_VGND_c_1154_n 0.0030414f $X=9.095 $Y=0.745 $X2=0 $Y2=0
cc_557 N_A2_N_M1020_g N_VGND_c_1154_n 0.0030414f $X=9.525 $Y=0.745 $X2=0 $Y2=0
cc_558 N_A2_N_M1001_g N_VGND_c_1155_n 0.00435814f $X=8.235 $Y=0.745 $X2=0 $Y2=0
cc_559 N_A2_N_M1016_g N_VGND_c_1155_n 0.0043484f $X=8.665 $Y=0.745 $X2=0 $Y2=0
cc_560 N_A2_N_M1018_g N_VGND_c_1155_n 0.0043393f $X=9.095 $Y=0.745 $X2=0 $Y2=0
cc_561 N_A2_N_M1020_g N_VGND_c_1155_n 0.004733f $X=9.525 $Y=0.745 $X2=0 $Y2=0
cc_562 N_A2_N_M1001_g N_A_1235_65#_c_1276_n 7.73317e-19 $X=8.235 $Y=0.745 $X2=0
+ $Y2=0
cc_563 N_A2_N_c_656_n N_A_1235_65#_c_1276_n 0.00660344f $X=8.763 $Y=1.382 $X2=0
+ $Y2=0
cc_564 N_A2_N_M1001_g N_A_1235_65#_c_1277_n 0.0117422f $X=8.235 $Y=0.745 $X2=0
+ $Y2=0
cc_565 N_A2_N_M1016_g N_A_1235_65#_c_1277_n 0.00871207f $X=8.665 $Y=0.745 $X2=0
+ $Y2=0
cc_566 N_A2_N_M1018_g N_A_1235_65#_c_1279_n 0.00861516f $X=9.095 $Y=0.745 $X2=0
+ $Y2=0
cc_567 N_A2_N_M1020_g N_A_1235_65#_c_1279_n 0.0127933f $X=9.525 $Y=0.745 $X2=0
+ $Y2=0
cc_568 N_A2_N_M1016_g N_A_1235_65#_c_1282_n 2.16803e-19 $X=8.665 $Y=0.745 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_735_n N_A_132_367#_M1009_s 0.00371719f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_570 N_VPWR_c_735_n N_A_132_367#_M1036_s 0.00281079f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_735_n N_A_132_367#_M1021_s 0.00223577f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_735_n N_A_132_367#_M1037_s 0.00223577f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_737_n N_A_132_367#_c_895_n 0.00122268f $X=0.37 $Y=1.98 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_753_n N_A_132_367#_c_922_n 0.0128073f $X=1.065 $Y=3.33 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_735_n N_A_132_367#_c_922_n 0.00768194f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_576 N_VPWR_M1012_d N_A_132_367#_c_905_n 0.00362265f $X=1.09 $Y=1.835 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_738_n N_A_132_367#_c_905_n 0.0166566f $X=1.23 $Y=2.815 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_735_n N_A_132_367#_c_905_n 0.011595f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_579 N_VPWR_c_747_n N_A_132_367#_c_927_n 0.014278f $X=3.745 $Y=3.33 $X2=0
+ $Y2=0
cc_580 N_VPWR_c_735_n N_A_132_367#_c_927_n 0.00815375f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_581 N_VPWR_c_747_n N_A_132_367#_c_911_n 0.100711f $X=3.745 $Y=3.33 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_735_n N_A_132_367#_c_911_n 0.0648018f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_735_n N_Y_M1005_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_584 N_VPWR_c_735_n N_Y_M1032_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_585 N_VPWR_c_735_n N_Y_M1002_d 0.00399203f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_586 N_VPWR_c_735_n N_Y_M1013_d 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_587 N_VPWR_c_749_n N_Y_c_993_n 0.0124525f $X=4.575 $Y=3.33 $X2=0 $Y2=0
cc_588 N_VPWR_c_735_n N_Y_c_993_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_589 N_VPWR_M1008_s N_Y_c_940_n 0.00176461f $X=4.6 $Y=1.835 $X2=0 $Y2=0
cc_590 N_VPWR_c_740_n N_Y_c_940_n 0.0170777f $X=4.74 $Y=2.21 $X2=0 $Y2=0
cc_591 N_VPWR_c_754_n N_Y_c_997_n 0.0124525f $X=5.435 $Y=3.33 $X2=0 $Y2=0
cc_592 N_VPWR_c_735_n N_Y_c_997_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_593 N_VPWR_M1038_d Y 0.00901569f $X=3.7 $Y=1.835 $X2=0 $Y2=0
cc_594 N_VPWR_c_739_n Y 0.0186197f $X=3.88 $Y=2.965 $X2=0 $Y2=0
cc_595 N_VPWR_c_747_n Y 0.0022051f $X=3.745 $Y=3.33 $X2=0 $Y2=0
cc_596 N_VPWR_c_749_n Y 0.00229776f $X=4.575 $Y=3.33 $X2=0 $Y2=0
cc_597 N_VPWR_c_735_n Y 0.0125386f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_598 N_VPWR_c_737_n N_A_35_65#_c_1022_n 7.2296e-19 $X=0.37 $Y=1.98 $X2=0 $Y2=0
cc_599 N_VPWR_c_737_n N_A_35_65#_c_1023_n 0.00484872f $X=0.37 $Y=1.98 $X2=0
+ $Y2=0
cc_600 N_A_132_367#_c_911_n N_Y_M1005_d 0.00337742f $X=3.41 $Y=2.915 $X2=0 $Y2=0
cc_601 N_A_132_367#_c_911_n N_Y_M1032_d 0.00337742f $X=3.41 $Y=2.915 $X2=0 $Y2=0
cc_602 N_A_132_367#_M1021_s Y 0.00347261f $X=2.41 $Y=1.835 $X2=0 $Y2=0
cc_603 N_A_132_367#_M1037_s Y 0.00353801f $X=3.27 $Y=1.835 $X2=0 $Y2=0
cc_604 N_A_132_367#_c_911_n Y 0.083757f $X=3.41 $Y=2.915 $X2=0 $Y2=0
cc_605 N_Y_c_937_n N_A_35_65#_M1023_d 0.00267852f $X=5.185 $Y=1.16 $X2=0 $Y2=0
cc_606 N_Y_c_936_n N_A_35_65#_c_1029_n 8.86177e-19 $X=4.08 $Y=1.775 $X2=0 $Y2=0
cc_607 N_Y_c_938_n N_A_35_65#_c_1029_n 0.0110535f $X=4.245 $Y=1.16 $X2=0 $Y2=0
cc_608 N_Y_c_965_n N_A_35_65#_c_1053_n 0.00732365f $X=4.33 $Y=0.7 $X2=0 $Y2=0
cc_609 N_Y_M1011_s N_A_35_65#_c_1030_n 0.00197722f $X=4.17 $Y=0.325 $X2=0 $Y2=0
cc_610 N_Y_c_965_n N_A_35_65#_c_1030_n 0.016037f $X=4.33 $Y=0.7 $X2=0 $Y2=0
cc_611 N_Y_c_937_n N_A_35_65#_c_1030_n 0.00280043f $X=5.185 $Y=1.16 $X2=0 $Y2=0
cc_612 N_Y_c_938_n N_A_35_65#_c_1030_n 0.00365354f $X=4.245 $Y=1.16 $X2=0 $Y2=0
cc_613 N_Y_c_937_n N_A_35_65#_c_1080_n 0.0207523f $X=5.185 $Y=1.16 $X2=0 $Y2=0
cc_614 N_Y_M1027_s N_A_35_65#_c_1032_n 0.00267852f $X=5.13 $Y=0.325 $X2=0 $Y2=0
cc_615 N_Y_c_937_n N_A_35_65#_c_1032_n 0.00280043f $X=5.185 $Y=1.16 $X2=0 $Y2=0
cc_616 N_Y_c_979_n N_A_35_65#_c_1032_n 0.0193433f $X=5.35 $Y=0.7 $X2=0 $Y2=0
cc_617 N_A_35_65#_c_1022_n N_VGND_M1017_s 0.00176773f $X=1.065 $Y=1.165
+ $X2=-0.19 $Y2=-0.245
cc_618 N_A_35_65#_c_1025_n N_VGND_M1034_s 0.00176773f $X=1.925 $Y=1.165 $X2=0
+ $Y2=0
cc_619 N_A_35_65#_c_1027_n N_VGND_M1015_s 0.00176773f $X=2.785 $Y=1.165 $X2=0
+ $Y2=0
cc_620 N_A_35_65#_c_1029_n N_VGND_M1030_s 0.00261503f $X=3.655 $Y=1.17 $X2=0
+ $Y2=0
cc_621 N_A_35_65#_c_1021_n N_VGND_c_1138_n 0.0222328f $X=0.3 $Y=0.47 $X2=0 $Y2=0
cc_622 N_A_35_65#_c_1022_n N_VGND_c_1138_n 0.0171443f $X=1.065 $Y=1.165 $X2=0
+ $Y2=0
cc_623 N_A_35_65#_c_1024_n N_VGND_c_1138_n 0.0232405f $X=1.16 $Y=0.47 $X2=0
+ $Y2=0
cc_624 N_A_35_65#_c_1024_n N_VGND_c_1139_n 0.0232405f $X=1.16 $Y=0.47 $X2=0
+ $Y2=0
cc_625 N_A_35_65#_c_1025_n N_VGND_c_1139_n 0.0171443f $X=1.925 $Y=1.165 $X2=0
+ $Y2=0
cc_626 N_A_35_65#_c_1026_n N_VGND_c_1139_n 0.0232405f $X=2.02 $Y=0.47 $X2=0
+ $Y2=0
cc_627 N_A_35_65#_c_1026_n N_VGND_c_1140_n 0.0232405f $X=2.02 $Y=0.47 $X2=0
+ $Y2=0
cc_628 N_A_35_65#_c_1027_n N_VGND_c_1140_n 0.0171443f $X=2.785 $Y=1.165 $X2=0
+ $Y2=0
cc_629 N_A_35_65#_c_1028_n N_VGND_c_1140_n 0.0232405f $X=2.88 $Y=0.47 $X2=0
+ $Y2=0
cc_630 N_A_35_65#_c_1028_n N_VGND_c_1141_n 0.0237205f $X=2.88 $Y=0.47 $X2=0
+ $Y2=0
cc_631 N_A_35_65#_c_1029_n N_VGND_c_1141_n 0.0218003f $X=3.655 $Y=1.17 $X2=0
+ $Y2=0
cc_632 N_A_35_65#_c_1031_n N_VGND_c_1141_n 0.00963725f $X=3.985 $Y=0.35 $X2=0
+ $Y2=0
cc_633 N_A_35_65#_c_1032_n N_VGND_c_1142_n 0.00126808f $X=5.685 $Y=0.35 $X2=0
+ $Y2=0
cc_634 N_A_35_65#_c_1024_n N_VGND_c_1145_n 0.0102275f $X=1.16 $Y=0.47 $X2=0
+ $Y2=0
cc_635 N_A_35_65#_c_1026_n N_VGND_c_1147_n 0.0102275f $X=2.02 $Y=0.47 $X2=0
+ $Y2=0
cc_636 N_A_35_65#_c_1028_n N_VGND_c_1149_n 0.0102275f $X=2.88 $Y=0.47 $X2=0
+ $Y2=0
cc_637 N_A_35_65#_c_1030_n N_VGND_c_1151_n 0.0409239f $X=4.675 $Y=0.35 $X2=0
+ $Y2=0
cc_638 N_A_35_65#_c_1031_n N_VGND_c_1151_n 0.0221146f $X=3.985 $Y=0.35 $X2=0
+ $Y2=0
cc_639 N_A_35_65#_c_1032_n N_VGND_c_1151_n 0.0579224f $X=5.685 $Y=0.35 $X2=0
+ $Y2=0
cc_640 N_A_35_65#_c_1037_n N_VGND_c_1151_n 0.0220373f $X=4.84 $Y=0.35 $X2=0
+ $Y2=0
cc_641 N_A_35_65#_c_1021_n N_VGND_c_1153_n 0.0134916f $X=0.3 $Y=0.47 $X2=0 $Y2=0
cc_642 N_A_35_65#_c_1021_n N_VGND_c_1155_n 0.0093995f $X=0.3 $Y=0.47 $X2=0 $Y2=0
cc_643 N_A_35_65#_c_1024_n N_VGND_c_1155_n 0.00712543f $X=1.16 $Y=0.47 $X2=0
+ $Y2=0
cc_644 N_A_35_65#_c_1026_n N_VGND_c_1155_n 0.00712543f $X=2.02 $Y=0.47 $X2=0
+ $Y2=0
cc_645 N_A_35_65#_c_1028_n N_VGND_c_1155_n 0.00712543f $X=2.88 $Y=0.47 $X2=0
+ $Y2=0
cc_646 N_A_35_65#_c_1030_n N_VGND_c_1155_n 0.0244057f $X=4.675 $Y=0.35 $X2=0
+ $Y2=0
cc_647 N_A_35_65#_c_1031_n N_VGND_c_1155_n 0.0126434f $X=3.985 $Y=0.35 $X2=0
+ $Y2=0
cc_648 N_A_35_65#_c_1032_n N_VGND_c_1155_n 0.0342072f $X=5.685 $Y=0.35 $X2=0
+ $Y2=0
cc_649 N_A_35_65#_c_1037_n N_VGND_c_1155_n 0.0126273f $X=4.84 $Y=0.35 $X2=0
+ $Y2=0
cc_650 N_A_35_65#_c_1033_n N_A_1235_65#_c_1273_n 0.0136671f $X=5.78 $Y=0.47
+ $X2=0 $Y2=0
cc_651 N_A_35_65#_c_1032_n N_A_1235_65#_c_1274_n 0.0104513f $X=5.685 $Y=0.35
+ $X2=0 $Y2=0
cc_652 N_A_35_65#_c_1033_n N_A_1235_65#_c_1274_n 0.0322343f $X=5.78 $Y=0.47
+ $X2=0 $Y2=0
cc_653 N_VGND_c_1142_n N_A_1235_65#_c_1274_n 0.0155838f $X=6.73 $Y=0.58 $X2=0
+ $Y2=0
cc_654 N_VGND_c_1151_n N_A_1235_65#_c_1274_n 0.0140356f $X=6.565 $Y=0 $X2=0
+ $Y2=0
cc_655 N_VGND_c_1155_n N_A_1235_65#_c_1274_n 0.00977851f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_656 N_VGND_M1003_s N_A_1235_65#_c_1299_n 0.00404696f $X=6.59 $Y=0.325 $X2=0
+ $Y2=0
cc_657 N_VGND_c_1142_n N_A_1235_65#_c_1299_n 0.0170777f $X=6.73 $Y=0.58 $X2=0
+ $Y2=0
cc_658 N_VGND_c_1142_n N_A_1235_65#_c_1275_n 0.0155484f $X=6.73 $Y=0.58 $X2=0
+ $Y2=0
cc_659 N_VGND_c_1143_n N_A_1235_65#_c_1275_n 0.0102275f $X=7.425 $Y=0 $X2=0
+ $Y2=0
cc_660 N_VGND_c_1144_n N_A_1235_65#_c_1275_n 0.0232405f $X=7.59 $Y=0.45 $X2=0
+ $Y2=0
cc_661 N_VGND_c_1155_n N_A_1235_65#_c_1275_n 0.00712543f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_662 N_VGND_M1024_s N_A_1235_65#_c_1276_n 0.00176461f $X=7.45 $Y=0.325 $X2=0
+ $Y2=0
cc_663 N_VGND_c_1144_n N_A_1235_65#_c_1276_n 0.0170777f $X=7.59 $Y=0.45 $X2=0
+ $Y2=0
cc_664 N_VGND_c_1154_n N_A_1235_65#_c_1277_n 0.0379195f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1155_n N_A_1235_65#_c_1277_n 0.0225412f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_666 N_VGND_c_1144_n N_A_1235_65#_c_1278_n 0.00915965f $X=7.59 $Y=0.45 $X2=0
+ $Y2=0
cc_667 N_VGND_c_1154_n N_A_1235_65#_c_1278_n 0.0128106f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_668 N_VGND_c_1155_n N_A_1235_65#_c_1278_n 0.0073517f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_669 N_VGND_c_1154_n N_A_1235_65#_c_1279_n 0.062494f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_670 N_VGND_c_1155_n N_A_1235_65#_c_1279_n 0.0367839f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_671 N_VGND_c_1154_n N_A_1235_65#_c_1282_n 0.0140519f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_672 N_VGND_c_1155_n N_A_1235_65#_c_1282_n 0.0083025f $X=9.84 $Y=0 $X2=0 $Y2=0
