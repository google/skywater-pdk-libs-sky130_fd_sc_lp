* File: sky130_fd_sc_lp__o21bai_2.pxi.spice
* Created: Fri Aug 28 11:06:43 2020
* 
x_PM_SKY130_FD_SC_LP__O21BAI_2%B1_N N_B1_N_c_79_n N_B1_N_M1013_g N_B1_N_c_80_n
+ N_B1_N_c_81_n N_B1_N_M1010_g B1_N B1_N N_B1_N_c_84_n N_B1_N_c_85_n
+ PM_SKY130_FD_SC_LP__O21BAI_2%B1_N
x_PM_SKY130_FD_SC_LP__O21BAI_2%A_100_367# N_A_100_367#_M1013_d
+ N_A_100_367#_M1010_s N_A_100_367#_c_108_n N_A_100_367#_M1006_g
+ N_A_100_367#_M1002_g N_A_100_367#_c_110_n N_A_100_367#_c_111_n
+ N_A_100_367#_M1012_g N_A_100_367#_M1009_g N_A_100_367#_c_113_n
+ N_A_100_367#_c_114_n N_A_100_367#_c_115_n N_A_100_367#_c_121_n
+ N_A_100_367#_c_116_n N_A_100_367#_c_117_n N_A_100_367#_c_118_n
+ PM_SKY130_FD_SC_LP__O21BAI_2%A_100_367#
x_PM_SKY130_FD_SC_LP__O21BAI_2%A1 N_A1_M1004_g N_A1_M1001_g N_A1_M1005_g
+ N_A1_M1003_g N_A1_c_186_n N_A1_c_179_n N_A1_c_180_n N_A1_c_181_n A1 A1 A1
+ N_A1_c_182_n N_A1_c_183_n A1 PM_SKY130_FD_SC_LP__O21BAI_2%A1
x_PM_SKY130_FD_SC_LP__O21BAI_2%A2 N_A2_M1000_g N_A2_M1008_g N_A2_M1007_g
+ N_A2_M1011_g A2 N_A2_c_263_n PM_SKY130_FD_SC_LP__O21BAI_2%A2
x_PM_SKY130_FD_SC_LP__O21BAI_2%VPWR N_VPWR_M1010_d N_VPWR_M1009_d N_VPWR_M1003_d
+ N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n VPWR
+ N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n
+ N_VPWR_c_312_n PM_SKY130_FD_SC_LP__O21BAI_2%VPWR
x_PM_SKY130_FD_SC_LP__O21BAI_2%Y N_Y_M1006_d N_Y_M1002_s N_Y_M1008_s N_Y_c_367_n
+ N_Y_c_390_n N_Y_c_369_n N_Y_c_370_n N_Y_c_365_n N_Y_c_364_n Y Y
+ PM_SKY130_FD_SC_LP__O21BAI_2%Y
x_PM_SKY130_FD_SC_LP__O21BAI_2%A_504_367# N_A_504_367#_M1001_s
+ N_A_504_367#_M1011_d N_A_504_367#_c_410_n N_A_504_367#_c_412_n
+ PM_SKY130_FD_SC_LP__O21BAI_2%A_504_367#
x_PM_SKY130_FD_SC_LP__O21BAI_2%VGND N_VGND_M1013_s N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n VGND
+ N_VGND_c_430_n N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n
+ N_VGND_c_435_n PM_SKY130_FD_SC_LP__O21BAI_2%VGND
x_PM_SKY130_FD_SC_LP__O21BAI_2%A_233_65# N_A_233_65#_M1006_s N_A_233_65#_M1012_s
+ N_A_233_65#_M1000_s N_A_233_65#_M1005_s N_A_233_65#_c_478_n
+ N_A_233_65#_c_479_n N_A_233_65#_c_480_n N_A_233_65#_c_481_n
+ N_A_233_65#_c_482_n N_A_233_65#_c_483_n N_A_233_65#_c_484_n
+ N_A_233_65#_c_485_n N_A_233_65#_c_486_n PM_SKY130_FD_SC_LP__O21BAI_2%A_233_65#
cc_1 VNB N_B1_N_c_79_n 0.0306189f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.36
cc_2 VNB N_B1_N_c_80_n 0.0243342f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.435
cc_3 VNB N_B1_N_c_81_n 0.0218451f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.435
cc_4 VNB N_B1_N_M1010_g 0.00868189f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.045
cc_5 VNB B1_N 0.041714f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B1_N_c_84_n 0.0235693f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_7 VNB N_B1_N_c_85_n 0.0241803f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=0.84
cc_8 VNB N_A_100_367#_c_108_n 0.0197518f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.435
cc_9 VNB N_A_100_367#_M1002_g 0.00293387f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_10 VNB N_A_100_367#_c_110_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_100_367#_c_111_n 0.0163952f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.005
cc_12 VNB N_A_100_367#_M1009_g 0.0115396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_100_367#_c_113_n 0.0052635f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.005
cc_14 VNB N_A_100_367#_c_114_n 0.0184957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_100_367#_c_115_n 0.0131082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_100_367#_c_116_n 0.00171733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_100_367#_c_117_n 0.00389865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_100_367#_c_118_n 0.0401613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1004_g 0.0204601f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_20 VNB N_A1_M1005_g 0.0261593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_179_n 0.00267096f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=0.84
cc_22 VNB N_A1_c_180_n 0.00849916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_181_n 0.0305833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_182_n 0.0245937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_183_n 0.00549405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_M1000_g 0.0206914f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_27 VNB N_A2_M1007_g 0.0192627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB A2 0.00155801f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_29 VNB N_A2_c_263_n 0.0313665f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_30 VNB N_VPWR_c_312_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_364_n 0.00493611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_426_n 0.0109343f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.045
cc_33 VNB N_VGND_c_427_n 0.0209936f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_34 VNB N_VGND_c_428_n 0.00458837f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.005
cc_35 VNB N_VGND_c_429_n 0.0023483f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_36 VNB N_VGND_c_430_n 0.0499053f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_37 VNB N_VGND_c_431_n 0.0161412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_432_n 0.0195242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_433_n 0.262082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_434_n 0.00586849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_435_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_233_65#_c_478_n 0.00941385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_233_65#_c_479_n 0.0047953f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_44 VNB N_A_233_65#_c_480_n 0.00453772f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_45 VNB N_A_233_65#_c_481_n 0.00463032f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.005
cc_46 VNB N_A_233_65#_c_482_n 0.00252946f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_47 VNB N_A_233_65#_c_483_n 0.00200294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_233_65#_c_484_n 0.0153442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_233_65#_c_485_n 0.0320667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_233_65#_c_486_n 0.00186402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_B1_N_M1010_g 0.0326067f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.045
cc_52 VPB N_A_100_367#_M1002_g 0.024065f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_53 VPB N_A_100_367#_M1009_g 0.020647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_100_367#_c_121_n 0.0209451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_100_367#_c_116_n 0.00346971f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A1_M1001_g 0.0183582f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.435
cc_57 VPB N_A1_M1003_g 0.0249715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A1_c_186_n 0.00136946f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.005
cc_59 VPB N_A1_c_181_n 0.00779349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A1_c_182_n 0.00638625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A1_c_183_n 0.00290651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A2_M1008_g 0.0183215f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.435
cc_63 VPB N_A2_M1011_g 0.0187184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB A2 0.00325047f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.005
cc_65 VPB N_A2_c_263_n 0.00469528f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_66 VPB N_VPWR_c_313_n 0.0446246f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_67 VPB N_VPWR_c_314_n 0.0027554f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.005
cc_68 VPB N_VPWR_c_315_n 0.013523f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_69 VPB N_VPWR_c_316_n 0.0557926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_317_n 0.0328515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_318_n 0.0141634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_319_n 0.0366357f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_320_n 0.0088221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_321_n 0.00516142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_312_n 0.0843754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_Y_c_365_n 8.40919e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_Y_c_364_n 0.00364643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 N_B1_N_M1010_g N_A_100_367#_M1002_g 0.00950166f $X=0.84 $Y=2.045 $X2=0
+ $Y2=0
cc_79 B1_N N_A_100_367#_c_114_n 0.0400018f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_B1_N_c_85_n N_A_100_367#_c_114_n 0.0175276f $X=0.362 $Y=0.84 $X2=0 $Y2=0
cc_81 N_B1_N_c_80_n N_A_100_367#_c_115_n 0.00302606f $X=0.765 $Y=1.435 $X2=0
+ $Y2=0
cc_82 N_B1_N_M1010_g N_A_100_367#_c_115_n 0.00407836f $X=0.84 $Y=2.045 $X2=0
+ $Y2=0
cc_83 N_B1_N_c_81_n N_A_100_367#_c_121_n 0.0053669f $X=0.55 $Y=1.435 $X2=0 $Y2=0
cc_84 N_B1_N_M1010_g N_A_100_367#_c_121_n 0.00878068f $X=0.84 $Y=2.045 $X2=0
+ $Y2=0
cc_85 N_B1_N_M1010_g N_A_100_367#_c_116_n 0.00575769f $X=0.84 $Y=2.045 $X2=0
+ $Y2=0
cc_86 N_B1_N_c_80_n N_A_100_367#_c_117_n 0.0161876f $X=0.765 $Y=1.435 $X2=0
+ $Y2=0
cc_87 N_B1_N_M1010_g N_A_100_367#_c_117_n 0.00558315f $X=0.84 $Y=2.045 $X2=0
+ $Y2=0
cc_88 B1_N N_A_100_367#_c_117_n 0.0123842f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_B1_N_c_79_n N_A_100_367#_c_118_n 0.00124058f $X=0.362 $Y=1.36 $X2=0
+ $Y2=0
cc_90 N_B1_N_c_80_n N_A_100_367#_c_118_n 0.0159229f $X=0.765 $Y=1.435 $X2=0
+ $Y2=0
cc_91 N_B1_N_M1010_g N_VPWR_c_313_n 0.0049024f $X=0.84 $Y=2.045 $X2=0 $Y2=0
cc_92 B1_N N_VGND_c_427_n 0.0257005f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_B1_N_c_84_n N_VGND_c_427_n 0.00158877f $X=0.34 $Y=1.005 $X2=0 $Y2=0
cc_94 N_B1_N_c_85_n N_VGND_c_427_n 0.0135644f $X=0.362 $Y=0.84 $X2=0 $Y2=0
cc_95 N_B1_N_c_85_n N_VGND_c_430_n 0.00425877f $X=0.362 $Y=0.84 $X2=0 $Y2=0
cc_96 B1_N N_VGND_c_433_n 0.00149795f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_97 N_B1_N_c_85_n N_VGND_c_433_n 0.00861707f $X=0.362 $Y=0.84 $X2=0 $Y2=0
cc_98 N_B1_N_c_85_n N_A_233_65#_c_480_n 0.00252129f $X=0.362 $Y=0.84 $X2=0 $Y2=0
cc_99 N_A_100_367#_c_111_n N_A1_M1004_g 0.0195151f $X=1.935 $Y=1.275 $X2=0 $Y2=0
cc_100 N_A_100_367#_M1009_g N_A1_M1001_g 0.0421636f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_101 N_A_100_367#_c_113_n N_A1_c_182_n 0.0174396f $X=1.935 $Y=1.35 $X2=0 $Y2=0
cc_102 N_A_100_367#_M1009_g N_A1_c_183_n 0.00526394f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_A_100_367#_M1002_g N_VPWR_c_313_n 0.00951624f $X=1.505 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_A_100_367#_c_115_n N_VPWR_c_313_n 0.0330105f $X=1.29 $Y=1.44 $X2=0
+ $Y2=0
cc_105 N_A_100_367#_c_121_n N_VPWR_c_313_n 0.0156867f $X=0.625 $Y=2.045 $X2=0
+ $Y2=0
cc_106 N_A_100_367#_c_118_n N_VPWR_c_313_n 0.0068226f $X=1.58 $Y=1.44 $X2=0
+ $Y2=0
cc_107 N_A_100_367#_M1002_g N_VPWR_c_314_n 5.3326e-19 $X=1.505 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_100_367#_M1009_g N_VPWR_c_314_n 0.00671141f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_A_100_367#_M1002_g N_VPWR_c_318_n 0.00585385f $X=1.505 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_100_367#_M1009_g N_VPWR_c_318_n 0.00391439f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_100_367#_M1002_g N_VPWR_c_312_n 0.0118084f $X=1.505 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_A_100_367#_M1009_g N_VPWR_c_312_n 0.00457021f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_100_367#_c_108_n N_Y_c_367_n 0.0045152f $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_114 N_A_100_367#_c_111_n N_Y_c_367_n 0.00429379f $X=1.935 $Y=1.275 $X2=0
+ $Y2=0
cc_115 N_A_100_367#_M1009_g N_Y_c_369_n 0.0199163f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_100_367#_c_108_n N_Y_c_370_n 0.00296571f $X=1.505 $Y=1.275 $X2=0
+ $Y2=0
cc_117 N_A_100_367#_c_111_n N_Y_c_370_n 0.00286104f $X=1.935 $Y=1.275 $X2=0
+ $Y2=0
cc_118 N_A_100_367#_M1002_g N_Y_c_365_n 4.976e-19 $X=1.505 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_100_367#_c_108_n N_Y_c_364_n 0.00244758f $X=1.505 $Y=1.275 $X2=0
+ $Y2=0
cc_120 N_A_100_367#_c_110_n N_Y_c_364_n 0.0146653f $X=1.86 $Y=1.35 $X2=0 $Y2=0
cc_121 N_A_100_367#_c_111_n N_Y_c_364_n 0.00129424f $X=1.935 $Y=1.275 $X2=0
+ $Y2=0
cc_122 N_A_100_367#_M1009_g N_Y_c_364_n 0.00352751f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_100_367#_c_115_n N_Y_c_364_n 0.0199243f $X=1.29 $Y=1.44 $X2=0 $Y2=0
cc_124 N_A_100_367#_c_118_n N_Y_c_364_n 0.00685975f $X=1.58 $Y=1.44 $X2=0 $Y2=0
cc_125 N_A_100_367#_c_111_n N_VGND_c_428_n 4.94886e-19 $X=1.935 $Y=1.275 $X2=0
+ $Y2=0
cc_126 N_A_100_367#_c_108_n N_VGND_c_430_n 0.00302501f $X=1.505 $Y=1.275 $X2=0
+ $Y2=0
cc_127 N_A_100_367#_c_111_n N_VGND_c_430_n 0.00302501f $X=1.935 $Y=1.275 $X2=0
+ $Y2=0
cc_128 N_A_100_367#_c_114_n N_VGND_c_430_n 0.0108042f $X=0.69 $Y=0.52 $X2=0
+ $Y2=0
cc_129 N_A_100_367#_c_108_n N_VGND_c_433_n 0.0048466f $X=1.505 $Y=1.275 $X2=0
+ $Y2=0
cc_130 N_A_100_367#_c_111_n N_VGND_c_433_n 0.00435646f $X=1.935 $Y=1.275 $X2=0
+ $Y2=0
cc_131 N_A_100_367#_c_114_n N_VGND_c_433_n 0.00950011f $X=0.69 $Y=0.52 $X2=0
+ $Y2=0
cc_132 N_A_100_367#_c_108_n N_A_233_65#_c_478_n 0.00352959f $X=1.505 $Y=1.275
+ $X2=0 $Y2=0
cc_133 N_A_100_367#_c_114_n N_A_233_65#_c_478_n 0.0440941f $X=0.69 $Y=0.52 $X2=0
+ $Y2=0
cc_134 N_A_100_367#_c_115_n N_A_233_65#_c_478_n 0.0205229f $X=1.29 $Y=1.44 $X2=0
+ $Y2=0
cc_135 N_A_100_367#_c_118_n N_A_233_65#_c_478_n 0.00636762f $X=1.58 $Y=1.44
+ $X2=0 $Y2=0
cc_136 N_A_100_367#_c_108_n N_A_233_65#_c_479_n 0.0125027f $X=1.505 $Y=1.275
+ $X2=0 $Y2=0
cc_137 N_A_100_367#_c_111_n N_A_233_65#_c_479_n 0.0118308f $X=1.935 $Y=1.275
+ $X2=0 $Y2=0
cc_138 N_A_100_367#_c_114_n N_A_233_65#_c_480_n 0.00440695f $X=0.69 $Y=0.52
+ $X2=0 $Y2=0
cc_139 N_A_100_367#_c_111_n N_A_233_65#_c_482_n 8.14086e-19 $X=1.935 $Y=1.275
+ $X2=0 $Y2=0
cc_140 N_A1_M1004_g N_A2_M1000_g 0.0237272f $X=2.365 $Y=0.745 $X2=0 $Y2=0
cc_141 N_A1_M1001_g N_A2_M1008_g 0.0544218f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_142 A1 N_A2_M1008_g 0.0110743f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_143 N_A1_c_183_n N_A2_M1008_g 0.0047115f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A1_M1005_g N_A2_M1007_g 0.024097f $X=3.735 $Y=0.745 $X2=0 $Y2=0
cc_145 N_A1_M1003_g N_A2_M1011_g 0.024097f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_146 A1 N_A2_M1011_g 0.0160255f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_147 N_A1_c_186_n A2 0.00812127f $X=3.605 $Y=1.92 $X2=0 $Y2=0
cc_148 N_A1_c_179_n A2 0.0186809f $X=3.695 $Y=1.535 $X2=0 $Y2=0
cc_149 N_A1_c_181_n A2 3.048e-19 $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_150 A1 A2 0.0369366f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_151 N_A1_c_182_n A2 8.84197e-19 $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_152 N_A1_c_183_n A2 0.0217414f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_153 N_A1_c_186_n N_A2_c_263_n 0.0043659f $X=3.605 $Y=1.92 $X2=0 $Y2=0
cc_154 N_A1_c_179_n N_A2_c_263_n 0.00174691f $X=3.695 $Y=1.535 $X2=0 $Y2=0
cc_155 N_A1_c_181_n N_A2_c_263_n 0.024097f $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_156 A1 N_A2_c_263_n 5.8554e-19 $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_157 N_A1_c_182_n N_A2_c_263_n 0.0208617f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A1_c_183_n N_A2_c_263_n 3.11791e-19 $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A1_c_183_n N_VPWR_M1009_d 0.004477f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A1_M1001_g N_VPWR_c_314_n 0.0047058f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A1_M1003_g N_VPWR_c_316_n 0.00858005f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A1_c_186_n N_VPWR_c_316_n 0.0043137f $X=3.605 $Y=1.92 $X2=0 $Y2=0
cc_163 N_A1_c_180_n N_VPWR_c_316_n 0.0101751f $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A1_c_181_n N_VPWR_c_316_n 0.00299509f $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A1_M1001_g N_VPWR_c_319_n 0.00422812f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A1_M1003_g N_VPWR_c_319_n 0.00547432f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A1_M1001_g N_VPWR_c_312_n 0.00610662f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A1_M1003_g N_VPWR_c_312_n 0.0108026f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_169 A1 N_Y_M1008_s 0.00334942f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_170 N_A1_M1001_g N_Y_c_369_n 0.0187059f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_171 A1 N_Y_c_369_n 0.0362406f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_172 N_A1_c_182_n N_Y_c_369_n 2.94749e-19 $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A1_c_183_n N_Y_c_369_n 0.0329808f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A1_M1004_g N_Y_c_364_n 3.16996e-19 $X=2.365 $Y=0.745 $X2=0 $Y2=0
cc_175 N_A1_c_182_n N_Y_c_364_n 3.99056e-19 $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A1_c_183_n N_Y_c_364_n 0.0344338f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_177 A1 N_A_504_367#_M1001_s 0.0056591f $X=3.515 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_178 N_A1_c_183_n N_A_504_367#_M1001_s 0.00168185f $X=2.415 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A1_c_186_n N_A_504_367#_M1011_d 0.00192365f $X=3.605 $Y=1.92 $X2=0
+ $Y2=0
cc_180 A1 N_A_504_367#_M1011_d 0.00245081f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_181 N_A1_M1001_g N_A_504_367#_c_410_n 0.00335806f $X=2.445 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A1_M1003_g N_A_504_367#_c_410_n 0.00320931f $X=3.735 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A1_M1003_g N_A_504_367#_c_412_n 0.00788554f $X=3.735 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A1_c_186_n N_A_504_367#_c_412_n 0.00989454f $X=3.605 $Y=1.92 $X2=0
+ $Y2=0
cc_185 A1 N_A_504_367#_c_412_n 0.00818555f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_186 N_A1_M1004_g N_VGND_c_428_n 0.00852655f $X=2.365 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A1_M1005_g N_VGND_c_429_n 0.0124972f $X=3.735 $Y=0.745 $X2=0 $Y2=0
cc_188 N_A1_M1004_g N_VGND_c_430_n 0.00481374f $X=2.365 $Y=0.745 $X2=0 $Y2=0
cc_189 N_A1_M1005_g N_VGND_c_432_n 0.00414769f $X=3.735 $Y=0.745 $X2=0 $Y2=0
cc_190 N_A1_M1004_g N_VGND_c_433_n 0.00912395f $X=2.365 $Y=0.745 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_VGND_c_433_n 0.00826786f $X=3.735 $Y=0.745 $X2=0 $Y2=0
cc_192 N_A1_M1004_g N_A_233_65#_c_479_n 5.98295e-19 $X=2.365 $Y=0.745 $X2=0
+ $Y2=0
cc_193 N_A1_M1004_g N_A_233_65#_c_481_n 0.0139576f $X=2.365 $Y=0.745 $X2=0 $Y2=0
cc_194 A1 N_A_233_65#_c_481_n 0.00536799f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_195 N_A1_c_182_n N_A_233_65#_c_481_n 0.00442212f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A1_c_183_n N_A_233_65#_c_481_n 0.0245374f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A1_c_182_n N_A_233_65#_c_482_n 3.84846e-19 $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_198 N_A1_c_183_n N_A_233_65#_c_482_n 0.0187018f $X=2.415 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A1_M1004_g N_A_233_65#_c_483_n 4.15588e-19 $X=2.365 $Y=0.745 $X2=0
+ $Y2=0
cc_200 N_A1_M1005_g N_A_233_65#_c_484_n 0.0140377f $X=3.735 $Y=0.745 $X2=0 $Y2=0
cc_201 N_A1_c_179_n N_A_233_65#_c_484_n 0.01494f $X=3.695 $Y=1.535 $X2=0 $Y2=0
cc_202 N_A1_c_180_n N_A_233_65#_c_484_n 0.0222364f $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_203 N_A1_c_181_n N_A_233_65#_c_484_n 0.00457279f $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_204 A1 N_A_233_65#_c_484_n 0.00375601f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_205 N_A1_M1005_g N_A_233_65#_c_485_n 0.00354659f $X=3.735 $Y=0.745 $X2=0
+ $Y2=0
cc_206 N_A2_M1008_g N_VPWR_c_319_n 0.00357877f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A2_M1011_g N_VPWR_c_319_n 0.00357842f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A2_M1008_g N_VPWR_c_312_n 0.00537654f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A2_M1011_g N_VPWR_c_312_n 0.00537652f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A2_M1008_g N_Y_c_369_n 0.0126738f $X=2.875 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A2_M1008_g N_A_504_367#_c_410_n 0.0105192f $X=2.875 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_A2_M1011_g N_A_504_367#_c_410_n 0.014133f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A2_M1008_g N_A_504_367#_c_412_n 8.1291e-19 $X=2.875 $Y=2.465 $X2=0
+ $Y2=0
cc_214 N_A2_M1011_g N_A_504_367#_c_412_n 0.00893026f $X=3.305 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_A2_M1000_g N_VGND_c_428_n 0.00492622f $X=2.875 $Y=0.745 $X2=0 $Y2=0
cc_216 N_A2_M1000_g N_VGND_c_429_n 6.06779e-19 $X=2.875 $Y=0.745 $X2=0 $Y2=0
cc_217 N_A2_M1007_g N_VGND_c_429_n 0.0102888f $X=3.305 $Y=0.745 $X2=0 $Y2=0
cc_218 N_A2_M1000_g N_VGND_c_431_n 0.0048189f $X=2.875 $Y=0.745 $X2=0 $Y2=0
cc_219 N_A2_M1007_g N_VGND_c_431_n 0.00414769f $X=3.305 $Y=0.745 $X2=0 $Y2=0
cc_220 N_A2_M1000_g N_VGND_c_433_n 0.0093244f $X=2.875 $Y=0.745 $X2=0 $Y2=0
cc_221 N_A2_M1007_g N_VGND_c_433_n 0.00787505f $X=3.305 $Y=0.745 $X2=0 $Y2=0
cc_222 N_A2_M1000_g N_A_233_65#_c_481_n 0.0122687f $X=2.875 $Y=0.745 $X2=0 $Y2=0
cc_223 A2 N_A_233_65#_c_481_n 0.00959498f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A2_M1000_g N_A_233_65#_c_483_n 0.0108894f $X=2.875 $Y=0.745 $X2=0 $Y2=0
cc_225 N_A2_M1007_g N_A_233_65#_c_483_n 8.32384e-19 $X=3.305 $Y=0.745 $X2=0
+ $Y2=0
cc_226 N_A2_M1007_g N_A_233_65#_c_484_n 0.0138139f $X=3.305 $Y=0.745 $X2=0 $Y2=0
cc_227 A2 N_A_233_65#_c_484_n 0.0115436f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_228 N_A2_M1000_g N_A_233_65#_c_486_n 0.00151304f $X=2.875 $Y=0.745 $X2=0
+ $Y2=0
cc_229 A2 N_A_233_65#_c_486_n 0.0209954f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_230 N_A2_c_263_n N_A_233_65#_c_486_n 0.00256759f $X=3.305 $Y=1.51 $X2=0 $Y2=0
cc_231 N_VPWR_c_312_n N_Y_M1002_s 0.00290842f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_232 N_VPWR_c_312_n N_Y_M1008_s 0.00225186f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_233 N_VPWR_c_318_n N_Y_c_390_n 0.0138717f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_234 N_VPWR_c_312_n N_Y_c_390_n 0.00886411f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_235 N_VPWR_M1009_d N_Y_c_369_n 0.00521003f $X=2.01 $Y=1.835 $X2=0 $Y2=0
cc_236 N_VPWR_c_314_n N_Y_c_369_n 0.0210565f $X=2.16 $Y=2.915 $X2=0 $Y2=0
cc_237 N_VPWR_c_318_n N_Y_c_369_n 0.00205271f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_238 N_VPWR_c_319_n N_Y_c_369_n 0.00215663f $X=3.865 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_312_n N_Y_c_369_n 0.0102509f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_240 N_VPWR_c_313_n N_Y_c_365_n 0.00158911f $X=1.055 $Y=1.98 $X2=0 $Y2=0
cc_241 N_VPWR_c_312_n Y 5.66896e-19 $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_312_n N_A_504_367#_M1001_s 0.00223577f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_243 N_VPWR_c_312_n N_A_504_367#_M1011_d 0.00223559f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_319_n N_A_504_367#_c_410_n 0.067688f $X=3.865 $Y=3.33 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_312_n N_A_504_367#_c_410_n 0.0435984f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_316_n N_A_233_65#_c_484_n 0.00505244f $X=3.95 $Y=1.98 $X2=0
+ $Y2=0
cc_247 N_Y_c_369_n N_A_504_367#_M1001_s 0.00354899f $X=3.09 $Y=2.455 $X2=-0.19
+ $Y2=-0.245
cc_248 N_Y_M1008_s N_A_504_367#_c_410_n 0.00342096f $X=2.95 $Y=1.835 $X2=0 $Y2=0
cc_249 N_Y_c_369_n N_A_504_367#_c_410_n 0.0355503f $X=3.09 $Y=2.455 $X2=0 $Y2=0
cc_250 N_Y_c_364_n N_A_233_65#_c_478_n 0.00114645f $X=1.72 $Y=1.815 $X2=0 $Y2=0
cc_251 N_Y_M1006_d N_A_233_65#_c_479_n 0.00176461f $X=1.58 $Y=0.325 $X2=0 $Y2=0
cc_252 N_Y_c_367_n N_A_233_65#_c_479_n 0.0159261f $X=1.72 $Y=0.68 $X2=0 $Y2=0
cc_253 N_Y_c_364_n N_A_233_65#_c_482_n 0.00637401f $X=1.72 $Y=1.815 $X2=0 $Y2=0
cc_254 N_VGND_c_428_n N_A_233_65#_c_479_n 0.00962579f $X=2.6 $Y=0.45 $X2=0 $Y2=0
cc_255 N_VGND_c_430_n N_A_233_65#_c_479_n 0.0578544f $X=2.435 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_433_n N_A_233_65#_c_479_n 0.0323448f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_430_n N_A_233_65#_c_480_n 0.0179217f $X=2.435 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_433_n N_A_233_65#_c_480_n 0.00971942f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_M1004_d N_A_233_65#_c_481_n 0.00261503f $X=2.44 $Y=0.325 $X2=0
+ $Y2=0
cc_260 N_VGND_c_428_n N_A_233_65#_c_481_n 0.0202768f $X=2.6 $Y=0.45 $X2=0 $Y2=0
cc_261 N_VGND_c_428_n N_A_233_65#_c_483_n 0.0227258f $X=2.6 $Y=0.45 $X2=0 $Y2=0
cc_262 N_VGND_c_429_n N_A_233_65#_c_483_n 0.0236466f $X=3.52 $Y=0.45 $X2=0 $Y2=0
cc_263 N_VGND_c_431_n N_A_233_65#_c_483_n 0.0134464f $X=3.355 $Y=0 $X2=0 $Y2=0
cc_264 N_VGND_c_433_n N_A_233_65#_c_483_n 0.00933346f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_M1007_d N_A_233_65#_c_484_n 0.00176461f $X=3.38 $Y=0.325 $X2=0
+ $Y2=0
cc_266 N_VGND_c_429_n N_A_233_65#_c_484_n 0.0170777f $X=3.52 $Y=0.45 $X2=0 $Y2=0
cc_267 N_VGND_c_429_n N_A_233_65#_c_485_n 0.0236597f $X=3.52 $Y=0.45 $X2=0 $Y2=0
cc_268 N_VGND_c_432_n N_A_233_65#_c_485_n 0.0151237f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_433_n N_A_233_65#_c_485_n 0.0105365f $X=4.08 $Y=0 $X2=0 $Y2=0
