# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xor2_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__xor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.370000 0.615000 3.920000 0.785000 ;
        RECT 0.370000 0.785000 0.540000 1.345000 ;
        RECT 0.370000 1.345000 0.845000 1.605000 ;
        RECT 0.675000 1.605000 0.845000 1.950000 ;
        RECT 0.675000 1.950000 2.335000 2.120000 ;
        RECT 1.595000 1.345000 2.335000 1.950000 ;
        RECT 3.740000 0.785000 3.920000 1.355000 ;
        RECT 3.740000 1.355000 4.070000 1.605000 ;
        RECT 3.900000 1.605000 4.070000 1.920000 ;
        RECT 3.900000 1.920000 5.725000 2.090000 ;
        RECT 5.395000 1.415000 5.725000 1.920000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.345000 1.425000 1.780000 ;
        RECT 4.285000 1.415000 4.955000 1.750000 ;
      LAYER mcon ;
        RECT 1.115000 1.580000 1.285000 1.750000 ;
        RECT 4.475000 1.580000 4.645000 1.750000 ;
      LAYER met1 ;
        RECT 1.055000 1.550000 1.345000 1.595000 ;
        RECT 1.055000 1.595000 4.705000 1.735000 ;
        RECT 1.055000 1.735000 1.345000 1.780000 ;
        RECT 4.415000 1.550000 4.705000 1.595000 ;
        RECT 4.415000 1.735000 4.705000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.844200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 0.955000 3.380000 1.160000 ;
        RECT 3.050000 1.840000 3.380000 2.260000 ;
        RECT 3.050000 2.260000 6.155000 2.430000 ;
        RECT 3.210000 1.160000 3.380000 1.840000 ;
        RECT 4.475000 0.595000 4.805000 0.810000 ;
        RECT 4.475000 0.810000 5.125000 1.075000 ;
        RECT 4.475000 1.075000 6.155000 1.245000 ;
        RECT 5.895000 1.245000 6.155000 2.260000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.240000 0.085000 ;
        RECT 0.195000  0.085000 0.525000 0.445000 ;
        RECT 1.230000  0.085000 1.560000 0.445000 ;
        RECT 2.480000  0.085000 2.810000 0.445000 ;
        RECT 3.535000  0.085000 3.865000 0.445000 ;
        RECT 5.795000  0.085000 6.125000 0.905000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.240000 3.415000 ;
        RECT 0.255000 1.820000 0.505000 2.290000 ;
        RECT 0.255000 2.290000 0.620000 3.245000 ;
        RECT 2.100000 2.630000 2.430000 3.245000 ;
        RECT 3.990000 2.940000 4.320000 3.245000 ;
        RECT 5.010000 2.940000 5.340000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.720000 0.955000 2.700000 1.175000 ;
      RECT 0.790000 2.290000 1.020000 2.800000 ;
      RECT 0.790000 2.800000 1.930000 3.075000 ;
      RECT 1.190000 2.290000 2.700000 2.460000 ;
      RECT 1.190000 2.460000 1.430000 2.630000 ;
      RECT 1.600000 2.630000 1.930000 2.800000 ;
      RECT 2.530000 1.175000 2.700000 1.330000 ;
      RECT 2.530000 1.330000 3.030000 1.605000 ;
      RECT 2.530000 1.605000 2.700000 2.290000 ;
      RECT 2.620000 2.630000 5.850000 2.770000 ;
      RECT 2.620000 2.770000 3.810000 3.075000 ;
      RECT 2.965000 2.600000 5.850000 2.630000 ;
      RECT 4.090000 0.255000 5.625000 0.425000 ;
      RECT 4.090000 0.425000 4.305000 1.185000 ;
      RECT 4.975000 0.425000 5.625000 0.640000 ;
      RECT 5.295000 0.640000 5.625000 0.905000 ;
  END
END sky130_fd_sc_lp__xor2_2
