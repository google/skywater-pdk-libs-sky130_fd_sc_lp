* NGSPICE file created from sky130_fd_sc_lp__and3_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and3_0 A B C VGND VNB VPB VPWR X
M1000 VPWR C a_68_65# VPB phighvt w=420000u l=150000u
+  ad=4.726e+11p pd=3.92e+06u as=2.289e+11p ps=2.77e+06u
M1001 VGND C a_229_65# VNB nshort w=420000u l=150000u
+  ad=3.465e+11p pd=2.49e+06u as=8.82e+10p ps=1.26e+06u
M1002 a_68_65# B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_229_65# B a_157_65# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 X a_68_65# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1005 a_157_65# A a_68_65# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.239e+11p ps=1.43e+06u
M1006 X a_68_65# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 VPWR A a_68_65# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

