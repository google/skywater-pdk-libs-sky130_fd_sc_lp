* File: sky130_fd_sc_lp__mux4_0.pxi.spice
* Created: Wed Sep  2 10:01:45 2020
* 
x_PM_SKY130_FD_SC_LP__MUX4_0%A2 N_A2_c_177_n N_A2_c_178_n N_A2_M1017_g
+ N_A2_M1015_g N_A2_c_176_n A2 N_A2_c_181_n PM_SKY130_FD_SC_LP__MUX4_0%A2
x_PM_SKY130_FD_SC_LP__MUX4_0%S0 N_S0_c_225_n N_S0_c_226_n N_S0_M1012_g
+ N_S0_M1014_g N_S0_c_228_n N_S0_c_229_n N_S0_c_242_n N_S0_M1020_g N_S0_M1007_g
+ N_S0_c_231_n N_S0_c_232_n N_S0_M1001_g N_S0_c_234_n N_S0_M1011_g N_S0_c_236_n
+ N_S0_c_237_n N_S0_c_245_n N_S0_c_246_n S0 S0 N_S0_c_239_n
+ PM_SKY130_FD_SC_LP__MUX4_0%S0
x_PM_SKY130_FD_SC_LP__MUX4_0%A_31_506# N_A_31_506#_M1014_s N_A_31_506#_M1012_s
+ N_A_31_506#_M1009_g N_A_31_506#_M1004_g N_A_31_506#_M1025_g
+ N_A_31_506#_M1003_g N_A_31_506#_c_388_n N_A_31_506#_c_389_n
+ N_A_31_506#_c_390_n N_A_31_506#_c_391_n N_A_31_506#_c_400_n
+ N_A_31_506#_c_401_n N_A_31_506#_c_392_n N_A_31_506#_c_393_n
+ N_A_31_506#_c_402_n N_A_31_506#_c_403_n N_A_31_506#_c_404_n
+ N_A_31_506#_c_405_n N_A_31_506#_c_406_n N_A_31_506#_c_407_n
+ N_A_31_506#_c_459_n N_A_31_506#_c_408_n N_A_31_506#_c_409_n
+ N_A_31_506#_c_410_n N_A_31_506#_c_394_n N_A_31_506#_c_411_n
+ N_A_31_506#_c_395_n N_A_31_506#_c_413_n PM_SKY130_FD_SC_LP__MUX4_0%A_31_506#
x_PM_SKY130_FD_SC_LP__MUX4_0%A3 N_A3_M1010_g N_A3_M1002_g A3 N_A3_c_583_n
+ PM_SKY130_FD_SC_LP__MUX4_0%A3
x_PM_SKY130_FD_SC_LP__MUX4_0%A1 N_A1_M1023_g N_A1_M1005_g N_A1_c_622_n A1 A1 A1
+ N_A1_c_624_n PM_SKY130_FD_SC_LP__MUX4_0%A1
x_PM_SKY130_FD_SC_LP__MUX4_0%A0 N_A0_c_673_n N_A0_M1013_g N_A0_c_675_n
+ N_A0_M1024_g A0 PM_SKY130_FD_SC_LP__MUX4_0%A0
x_PM_SKY130_FD_SC_LP__MUX4_0%A_1029_37# N_A_1029_37#_M1021_s
+ N_A_1029_37#_M1022_s N_A_1029_37#_M1016_g N_A_1029_37#_M1000_g
+ N_A_1029_37#_c_719_n N_A_1029_37#_c_720_n N_A_1029_37#_c_711_n
+ N_A_1029_37#_c_712_n N_A_1029_37#_c_713_n N_A_1029_37#_c_714_n
+ N_A_1029_37#_c_723_n N_A_1029_37#_c_724_n N_A_1029_37#_c_715_n
+ N_A_1029_37#_c_716_n N_A_1029_37#_c_717_n
+ PM_SKY130_FD_SC_LP__MUX4_0%A_1029_37#
x_PM_SKY130_FD_SC_LP__MUX4_0%S1 N_S1_M1018_g N_S1_c_803_n N_S1_c_804_n
+ N_S1_c_805_n N_S1_M1006_g N_S1_c_806_n N_S1_M1022_g N_S1_M1021_g N_S1_c_808_n
+ N_S1_c_809_n N_S1_c_814_n S1 S1 S1 N_S1_c_811_n PM_SKY130_FD_SC_LP__MUX4_0%S1
x_PM_SKY130_FD_SC_LP__MUX4_0%A_1075_493# N_A_1075_493#_M1016_d
+ N_A_1075_493#_M1018_d N_A_1075_493#_c_904_n N_A_1075_493#_M1008_g
+ N_A_1075_493#_M1019_g N_A_1075_493#_c_900_n N_A_1075_493#_c_901_n
+ N_A_1075_493#_c_902_n N_A_1075_493#_c_907_n N_A_1075_493#_c_903_n
+ N_A_1075_493#_c_909_n N_A_1075_493#_c_914_n N_A_1075_493#_c_910_n
+ N_A_1075_493#_c_911_n N_A_1075_493#_c_912_n
+ PM_SKY130_FD_SC_LP__MUX4_0%A_1075_493#
x_PM_SKY130_FD_SC_LP__MUX4_0%VPWR N_VPWR_M1012_d N_VPWR_M1010_d N_VPWR_M1013_d
+ N_VPWR_M1022_d N_VPWR_c_976_n N_VPWR_c_977_n N_VPWR_c_978_n N_VPWR_c_979_n
+ N_VPWR_c_980_n N_VPWR_c_981_n N_VPWR_c_982_n N_VPWR_c_983_n N_VPWR_c_984_n
+ VPWR N_VPWR_c_985_n N_VPWR_c_986_n N_VPWR_c_987_n N_VPWR_c_975_n
+ N_VPWR_c_989_n N_VPWR_c_990_n N_VPWR_c_991_n PM_SKY130_FD_SC_LP__MUX4_0%VPWR
x_PM_SKY130_FD_SC_LP__MUX4_0%A_294_506# N_A_294_506#_M1009_d
+ N_A_294_506#_M1006_d N_A_294_506#_M1020_d N_A_294_506#_M1000_d
+ N_A_294_506#_c_1073_n N_A_294_506#_c_1065_n N_A_294_506#_c_1066_n
+ N_A_294_506#_c_1075_n N_A_294_506#_c_1067_n N_A_294_506#_c_1068_n
+ N_A_294_506#_c_1069_n N_A_294_506#_c_1070_n N_A_294_506#_c_1071_n
+ N_A_294_506#_c_1072_n PM_SKY130_FD_SC_LP__MUX4_0%A_294_506#
x_PM_SKY130_FD_SC_LP__MUX4_0%A_685_504# N_A_685_504#_M1001_d
+ N_A_685_504#_M1016_s N_A_685_504#_M1025_d N_A_685_504#_M1018_s
+ N_A_685_504#_c_1196_n N_A_685_504#_c_1185_n N_A_685_504#_c_1188_n
+ N_A_685_504#_c_1189_n N_A_685_504#_c_1186_n N_A_685_504#_c_1191_n
+ N_A_685_504#_c_1192_n N_A_685_504#_c_1187_n N_A_685_504#_c_1193_n
+ N_A_685_504#_c_1204_n N_A_685_504#_c_1205_n N_A_685_504#_c_1194_n
+ N_A_685_504#_c_1195_n PM_SKY130_FD_SC_LP__MUX4_0%A_685_504#
x_PM_SKY130_FD_SC_LP__MUX4_0%X N_X_M1008_d N_X_M1019_d X X X X X N_X_c_1275_n
+ PM_SKY130_FD_SC_LP__MUX4_0%X
x_PM_SKY130_FD_SC_LP__MUX4_0%VGND N_VGND_M1014_d N_VGND_M1002_d N_VGND_M1024_d
+ N_VGND_M1021_d N_VGND_c_1293_n N_VGND_c_1294_n N_VGND_c_1295_n N_VGND_c_1296_n
+ N_VGND_c_1297_n N_VGND_c_1298_n VGND N_VGND_c_1299_n N_VGND_c_1300_n
+ N_VGND_c_1301_n N_VGND_c_1302_n N_VGND_c_1303_n N_VGND_c_1304_n
+ N_VGND_c_1305_n N_VGND_c_1306_n PM_SKY130_FD_SC_LP__MUX4_0%VGND
cc_1 VNB N_A2_M1015_g 0.0339944f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=0.805
cc_2 VNB N_A2_c_176_n 0.0136574f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.625
cc_3 VNB N_S0_c_225_n 0.0156876f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.915
cc_4 VNB N_S0_c_226_n 0.00812063f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.305
cc_5 VNB N_S0_M1014_g 0.039067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_S0_c_228_n 0.0842518f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.625
cc_7 VNB N_S0_c_229_n 0.0126405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_S0_M1007_g 0.0363099f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.08
cc_9 VNB N_S0_c_231_n 0.0965572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_S0_c_232_n 0.0219236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_S0_M1001_g 0.0252406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_S0_c_234_n 0.0214507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_S0_M1011_g 0.00640928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_S0_c_236_n 0.0309671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_S0_c_237_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB S0 0.00279203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_S0_c_239_n 0.00279642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_31_506#_M1009_g 0.0266615f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=0.805
cc_19 VNB N_A_31_506#_M1003_g 0.027515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_31_506#_c_388_n 0.0621973f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.06
cc_21 VNB N_A_31_506#_c_389_n 0.00962308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_31_506#_c_390_n 0.0760615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_31_506#_c_391_n 0.0217244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_31_506#_c_392_n 0.0155589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_31_506#_c_393_n 0.0236495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_31_506#_c_394_n 0.0245162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_31_506#_c_395_n 0.0379978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A3_M1002_g 0.0452719f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.55
cc_29 VNB N_A1_M1005_g 0.017717f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.55
cc_30 VNB N_A1_c_622_n 0.0219375f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.625
cc_31 VNB A1 0.0103824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_c_624_n 0.0150466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A0_c_673_n 0.043574f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.7
cc_34 VNB N_A0_M1013_g 0.0019612f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.305
cc_35 VNB N_A0_c_675_n 0.0150618f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.74
cc_36 VNB A0 0.00452091f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=0.805
cc_37 VNB N_A_1029_37#_c_711_n 0.041074f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.08
cc_38 VNB N_A_1029_37#_c_712_n 0.0138134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1029_37#_c_713_n 0.0144789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1029_37#_c_714_n 9.79655e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1029_37#_c_715_n 0.0181467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1029_37#_c_716_n 0.00433158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1029_37#_c_717_n 0.0161977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_S1_M1018_g 0.00531877f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.305
cc_45 VNB N_S1_c_803_n 0.0220861f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.74
cc_46 VNB N_S1_c_804_n 0.00774051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_S1_c_805_n 0.0190363f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.55
cc_48 VNB N_S1_c_806_n 0.0430301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_S1_M1021_g 0.0425416f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.08
cc_50 VNB N_S1_c_808_n 0.0228164f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.06
cc_51 VNB N_S1_c_809_n 0.00966725f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.06
cc_52 VNB S1 0.0120867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_S1_c_811_n 0.0235226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1075_493#_c_900_n 0.0194906f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.08
cc_55 VNB N_A_1075_493#_c_901_n 0.0125674f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.08
cc_56 VNB N_A_1075_493#_c_902_n 0.0463276f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.06
cc_57 VNB N_A_1075_493#_c_903_n 0.00707647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VPWR_c_975_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_294_506#_c_1065_n 0.00643181f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=2.08
cc_60 VNB N_A_294_506#_c_1066_n 0.00262675f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=2.06
cc_61 VNB N_A_294_506#_c_1067_n 0.0026682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_294_506#_c_1068_n 0.00632042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_294_506#_c_1069_n 0.00390733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_294_506#_c_1070_n 0.00186621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_294_506#_c_1071_n 0.00346137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_294_506#_c_1072_n 0.00124729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_685_504#_c_1185_n 0.00586716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_685_504#_c_1186_n 0.00627007f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=2.08
cc_69 VNB N_A_685_504#_c_1187_n 0.0129428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_X_c_1275_n 0.0560176f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.08
cc_71 VNB N_VGND_c_1293_n 0.00831555f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_72 VNB N_VGND_c_1294_n 0.0105447f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.08
cc_73 VNB N_VGND_c_1295_n 0.0102607f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.06
cc_74 VNB N_VGND_c_1296_n 0.00519343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1297_n 0.0411444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1298_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1299_n 0.02844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1300_n 0.038647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1301_n 0.0532227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1302_n 0.0174529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1303_n 0.402653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1304_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1305_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1306_n 0.00487954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VPB N_A2_c_177_n 0.0130408f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=1.915
cc_86 VPB N_A2_c_178_n 0.0323752f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.305
cc_87 VPB N_A2_M1017_g 0.0213263f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.74
cc_88 VPB N_A2_c_176_n 0.00957538f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.625
cc_89 VPB N_A2_c_181_n 0.00500586f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.08
cc_90 VPB N_S0_c_226_n 0.0218972f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.305
cc_91 VPB N_S0_M1012_g 0.0485979f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.74
cc_92 VPB N_S0_c_242_n 0.0395088f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.625
cc_93 VPB N_S0_M1020_g 0.023109f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_94 VPB N_S0_M1011_g 0.0560055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_S0_c_245_n 0.00382616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_S0_c_246_n 0.00432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB S0 0.0039445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_S0_c_239_n 0.00304621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_31_506#_M1004_g 0.0525908f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.625
cc_100 VPB N_A_31_506#_M1025_g 0.0186107f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.08
cc_101 VPB N_A_31_506#_c_390_n 0.0124881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_31_506#_c_391_n 0.0342436f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_31_506#_c_400_n 0.0148572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_31_506#_c_401_n 0.0112961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_31_506#_c_402_n 0.00909221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_31_506#_c_403_n 0.00201781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_31_506#_c_404_n 0.0057976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_31_506#_c_405_n 8.37112e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_31_506#_c_406_n 0.0172177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_31_506#_c_407_n 0.00152567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_31_506#_c_408_n 0.0335548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_31_506#_c_409_n 0.00426898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_31_506#_c_410_n 0.0131502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_31_506#_c_411_n 0.0116996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_31_506#_c_395_n 0.0168589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_31_506#_c_413_n 0.0357372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A3_M1010_g 0.0252541f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.305
cc_118 VPB N_A3_M1002_g 0.0113023f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.55
cc_119 VPB A3 0.00609018f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=0.805
cc_120 VPB N_A3_c_583_n 0.0314221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A1_M1023_g 0.0353269f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.305
cc_122 VPB N_A1_c_622_n 0.0331511f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=1.625
cc_123 VPB A1 0.00791598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A0_M1013_g 0.0588845f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.305
cc_125 VPB N_A_1029_37#_M1000_g 0.0451967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_1029_37#_c_719_n 0.0167535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_1029_37#_c_720_n 0.00773947f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_128 VPB N_A_1029_37#_c_713_n 0.0299708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_1029_37#_c_714_n 0.00161376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_1029_37#_c_723_n 0.00408702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_1029_37#_c_724_n 0.00295844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_S1_M1018_g 0.0569519f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.305
cc_133 VPB N_S1_M1022_g 0.0224845f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_S1_c_814_n 0.0154369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB S1 0.00646976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_1075_493#_c_904_n 0.0425235f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=1.55
cc_137 VPB N_A_1075_493#_M1019_g 0.0164086f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_138 VPB N_A_1075_493#_c_902_n 0.00612751f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.06
cc_139 VPB N_A_1075_493#_c_907_n 0.012762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_1075_493#_c_903_n 0.0144267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_1075_493#_c_909_n 0.00530113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_1075_493#_c_910_n 0.00325071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1075_493#_c_911_n 0.0198259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_1075_493#_c_912_n 0.0440375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_976_n 0.0100484f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_146 VPB N_VPWR_c_977_n 0.00653909f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.08
cc_147 VPB N_VPWR_c_978_n 0.0135173f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.06
cc_148 VPB N_VPWR_c_979_n 0.0575999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_980_n 0.00460451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_981_n 0.00308069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_982_n 0.0157896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_983_n 0.0417238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_984_n 0.00474858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_985_n 0.0195023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_986_n 0.0408814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_987_n 0.0194843f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_975_n 0.113229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_989_n 0.00632327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_990_n 0.00628367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_991_n 0.00343303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_294_506#_c_1073_n 0.0126211f $X=-0.19 $Y=1.655 $X2=1.275
+ $Y2=1.625
cc_162 VPB N_A_294_506#_c_1065_n 0.00642795f $X=-0.19 $Y=1.655 $X2=0.945
+ $Y2=2.08
cc_163 VPB N_A_294_506#_c_1075_n 0.0107537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_294_506#_c_1067_n 0.00644126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_685_504#_c_1188_n 0.019981f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.08
cc_166 VPB N_A_685_504#_c_1189_n 0.00226814f $X=-0.19 $Y=1.655 $X2=0.945
+ $Y2=2.08
cc_167 VPB N_A_685_504#_c_1186_n 0.00562483f $X=-0.19 $Y=1.655 $X2=0.945
+ $Y2=2.08
cc_168 VPB N_A_685_504#_c_1191_n 6.95955e-19 $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.06
cc_169 VPB N_A_685_504#_c_1192_n 0.00501346f $X=-0.19 $Y=1.655 $X2=0.945
+ $Y2=2.06
cc_170 VPB N_A_685_504#_c_1193_n 0.00500269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_685_504#_c_1194_n 0.00288277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_685_504#_c_1195_n 0.001838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_X_c_1275_n 0.0451096f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.08
cc_174 N_A2_M1015_g N_S0_c_225_n 0.0047528f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_175 N_A2_c_177_n N_S0_c_226_n 0.00684995f $X=1.035 $Y=1.915 $X2=0 $Y2=0
cc_176 N_A2_c_176_n N_S0_c_226_n 0.00850429f $X=1.275 $Y=1.625 $X2=0 $Y2=0
cc_177 N_A2_c_181_n N_S0_c_226_n 9.34892e-19 $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_178 N_A2_c_178_n N_S0_M1012_g 0.0236336f $X=1.035 $Y=2.305 $X2=0 $Y2=0
cc_179 N_A2_M1017_g N_S0_M1012_g 0.0156353f $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_180 N_A2_c_181_n N_S0_M1012_g 0.00610174f $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_181 N_A2_M1015_g N_S0_M1014_g 0.0244045f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_182 N_A2_M1015_g N_S0_c_228_n 0.0103107f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_183 N_A2_c_178_n N_S0_c_242_n 0.0387039f $X=1.035 $Y=2.305 $X2=0 $Y2=0
cc_184 N_A2_c_176_n N_S0_c_242_n 6.88446e-19 $X=1.275 $Y=1.625 $X2=0 $Y2=0
cc_185 N_A2_c_181_n N_S0_c_242_n 2.80558e-19 $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_186 N_A2_M1017_g N_S0_M1020_g 0.0268726f $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_187 N_A2_c_178_n N_S0_c_236_n 0.00193743f $X=1.035 $Y=2.305 $X2=0 $Y2=0
cc_188 N_A2_c_177_n N_S0_c_245_n 0.00581044f $X=1.035 $Y=1.915 $X2=0 $Y2=0
cc_189 N_A2_c_181_n N_S0_c_245_n 6.78097e-19 $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_190 N_A2_c_178_n N_S0_c_246_n 8.72387e-19 $X=1.035 $Y=2.305 $X2=0 $Y2=0
cc_191 N_A2_c_181_n N_S0_c_246_n 0.0199842f $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_192 N_A2_c_177_n S0 0.00146679f $X=1.035 $Y=1.915 $X2=0 $Y2=0
cc_193 N_A2_M1015_g S0 0.0074162f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_194 N_A2_c_176_n S0 0.0111487f $X=1.275 $Y=1.625 $X2=0 $Y2=0
cc_195 N_A2_c_181_n S0 8.99751e-19 $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_196 N_A2_c_177_n N_S0_c_239_n 0.00350356f $X=1.035 $Y=1.915 $X2=0 $Y2=0
cc_197 N_A2_c_178_n N_S0_c_239_n 0.00239663f $X=1.035 $Y=2.305 $X2=0 $Y2=0
cc_198 N_A2_c_176_n N_S0_c_239_n 0.00593249f $X=1.275 $Y=1.625 $X2=0 $Y2=0
cc_199 N_A2_c_181_n N_S0_c_239_n 0.0433078f $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_200 N_A2_M1015_g N_A_31_506#_M1009_g 0.0374789f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_201 N_A2_c_181_n N_A_31_506#_c_391_n 0.0152732f $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_202 N_A2_M1017_g N_A_31_506#_c_400_n 6.12171e-19 $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_203 N_A2_c_178_n N_A_31_506#_c_401_n 0.00438639f $X=1.035 $Y=2.305 $X2=0
+ $Y2=0
cc_204 N_A2_M1017_g N_A_31_506#_c_401_n 0.0113969f $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_205 N_A2_c_176_n N_A_31_506#_c_401_n 0.00102128f $X=1.275 $Y=1.625 $X2=0
+ $Y2=0
cc_206 N_A2_c_181_n N_A_31_506#_c_401_n 0.0415361f $X=0.945 $Y=2.08 $X2=0 $Y2=0
cc_207 N_A2_M1015_g N_A_31_506#_c_393_n 0.0178028f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_208 N_A2_c_176_n N_A_31_506#_c_393_n 0.00112622f $X=1.275 $Y=1.625 $X2=0
+ $Y2=0
cc_209 N_A2_M1017_g N_A_31_506#_c_403_n 0.00115544f $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_210 N_A2_M1015_g N_A_31_506#_c_404_n 6.52111e-19 $X=1.275 $Y=0.805 $X2=0
+ $Y2=0
cc_211 N_A2_c_176_n N_A_31_506#_c_395_n 0.0374789f $X=1.275 $Y=1.625 $X2=0 $Y2=0
cc_212 N_A2_M1017_g N_VPWR_c_976_n 0.00139063f $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_213 N_A2_M1017_g N_VPWR_c_983_n 0.00570944f $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_214 N_A2_M1017_g N_VPWR_c_975_n 0.00542671f $X=1.035 $Y=2.74 $X2=0 $Y2=0
cc_215 N_A2_M1015_g N_VGND_c_1293_n 0.00917365f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_216 N_A2_M1015_g N_VGND_c_1303_n 7.88961e-19 $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_217 N_S0_c_228_n N_A_31_506#_M1009_g 0.0104164f $X=2.06 $Y=0.18 $X2=0 $Y2=0
cc_218 N_S0_M1007_g N_A_31_506#_M1009_g 0.015726f $X=2.135 $Y=0.805 $X2=0 $Y2=0
cc_219 N_S0_c_242_n N_A_31_506#_M1004_g 0.0146261f $X=1.395 $Y=2.305 $X2=0 $Y2=0
cc_220 N_S0_M1020_g N_A_31_506#_M1004_g 0.0151015f $X=1.395 $Y=2.74 $X2=0 $Y2=0
cc_221 N_S0_c_245_n N_A_31_506#_M1004_g 0.0026851f $X=1.375 $Y=1.94 $X2=0 $Y2=0
cc_222 N_S0_c_246_n N_A_31_506#_M1004_g 8.54127e-19 $X=1.515 $Y=2.105 $X2=0
+ $Y2=0
cc_223 S0 N_A_31_506#_M1004_g 0.00109093f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_224 N_S0_M1011_g N_A_31_506#_M1025_g 0.0103997f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_225 N_S0_c_232_n N_A_31_506#_M1003_g 0.0010151f $X=3.495 $Y=1.125 $X2=0 $Y2=0
cc_226 N_S0_M1001_g N_A_31_506#_M1003_g 0.0157854f $X=3.495 $Y=0.805 $X2=0 $Y2=0
cc_227 N_S0_c_234_n N_A_31_506#_M1003_g 0.00658315f $X=3.815 $Y=1.46 $X2=0 $Y2=0
cc_228 N_S0_c_231_n N_A_31_506#_c_389_n 0.0157854f $X=3.42 $Y=0.18 $X2=0 $Y2=0
cc_229 N_S0_M1012_g N_A_31_506#_c_391_n 0.0122952f $X=0.495 $Y=2.74 $X2=0 $Y2=0
cc_230 N_S0_c_236_n N_A_31_506#_c_391_n 0.0226741f $X=0.845 $Y=1.265 $X2=0 $Y2=0
cc_231 N_S0_c_239_n N_A_31_506#_c_391_n 0.03075f $X=1.098 $Y=1.567 $X2=0 $Y2=0
cc_232 N_S0_M1012_g N_A_31_506#_c_400_n 0.0060561f $X=0.495 $Y=2.74 $X2=0 $Y2=0
cc_233 N_S0_M1012_g N_A_31_506#_c_401_n 0.0107531f $X=0.495 $Y=2.74 $X2=0 $Y2=0
cc_234 N_S0_M1020_g N_A_31_506#_c_401_n 0.00424845f $X=1.395 $Y=2.74 $X2=0 $Y2=0
cc_235 N_S0_c_246_n N_A_31_506#_c_401_n 0.00130641f $X=1.515 $Y=2.105 $X2=0
+ $Y2=0
cc_236 S0 N_A_31_506#_c_401_n 0.006603f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_237 N_S0_c_239_n N_A_31_506#_c_401_n 0.00203845f $X=1.098 $Y=1.567 $X2=0
+ $Y2=0
cc_238 N_S0_M1014_g N_A_31_506#_c_392_n 6.81439e-19 $X=0.845 $Y=0.805 $X2=0
+ $Y2=0
cc_239 N_S0_c_236_n N_A_31_506#_c_392_n 0.00126872f $X=0.845 $Y=1.265 $X2=0
+ $Y2=0
cc_240 N_S0_M1014_g N_A_31_506#_c_393_n 0.0134547f $X=0.845 $Y=0.805 $X2=0 $Y2=0
cc_241 N_S0_c_242_n N_A_31_506#_c_393_n 0.00146218f $X=1.395 $Y=2.305 $X2=0
+ $Y2=0
cc_242 N_S0_c_236_n N_A_31_506#_c_393_n 0.00288549f $X=0.845 $Y=1.265 $X2=0
+ $Y2=0
cc_243 N_S0_c_246_n N_A_31_506#_c_393_n 0.00421786f $X=1.515 $Y=2.105 $X2=0
+ $Y2=0
cc_244 S0 N_A_31_506#_c_393_n 0.0221564f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_245 N_S0_c_242_n N_A_31_506#_c_402_n 0.00167925f $X=1.395 $Y=2.305 $X2=0
+ $Y2=0
cc_246 N_S0_M1020_g N_A_31_506#_c_402_n 0.0137074f $X=1.395 $Y=2.74 $X2=0 $Y2=0
cc_247 N_S0_c_246_n N_A_31_506#_c_404_n 0.00272701f $X=1.515 $Y=2.105 $X2=0
+ $Y2=0
cc_248 S0 N_A_31_506#_c_404_n 0.0175154f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_249 N_S0_M1011_g N_A_31_506#_c_406_n 5.60682e-19 $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_250 N_S0_M1011_g N_A_31_506#_c_459_n 7.85405e-19 $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_251 N_S0_c_232_n N_A_31_506#_c_408_n 0.00305606f $X=3.495 $Y=1.125 $X2=0
+ $Y2=0
cc_252 N_S0_M1011_g N_A_31_506#_c_408_n 0.0212887f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_253 N_S0_c_232_n N_A_31_506#_c_409_n 3.09793e-19 $X=3.495 $Y=1.125 $X2=0
+ $Y2=0
cc_254 N_S0_c_232_n N_A_31_506#_c_410_n 5.06683e-19 $X=3.495 $Y=1.125 $X2=0
+ $Y2=0
cc_255 N_S0_c_234_n N_A_31_506#_c_410_n 0.00362184f $X=3.815 $Y=1.46 $X2=0 $Y2=0
cc_256 N_S0_M1011_g N_A_31_506#_c_410_n 0.0144258f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_257 N_S0_M1014_g N_A_31_506#_c_394_n 4.14804e-19 $X=0.845 $Y=0.805 $X2=0
+ $Y2=0
cc_258 N_S0_c_236_n N_A_31_506#_c_394_n 0.0135813f $X=0.845 $Y=1.265 $X2=0 $Y2=0
cc_259 N_S0_c_239_n N_A_31_506#_c_394_n 0.0476592f $X=1.098 $Y=1.567 $X2=0 $Y2=0
cc_260 N_S0_c_226_n N_A_31_506#_c_411_n 0.00105278f $X=0.495 $Y=1.915 $X2=0
+ $Y2=0
cc_261 N_S0_M1012_g N_A_31_506#_c_411_n 0.00502934f $X=0.495 $Y=2.74 $X2=0 $Y2=0
cc_262 N_S0_c_242_n N_A_31_506#_c_395_n 0.00635351f $X=1.395 $Y=2.305 $X2=0
+ $Y2=0
cc_263 N_S0_M1007_g N_A_31_506#_c_395_n 0.00457864f $X=2.135 $Y=0.805 $X2=0
+ $Y2=0
cc_264 N_S0_c_246_n N_A_31_506#_c_395_n 4.22353e-19 $X=1.515 $Y=2.105 $X2=0
+ $Y2=0
cc_265 S0 N_A_31_506#_c_395_n 0.00154067f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_266 N_S0_M1007_g N_A3_M1002_g 0.0418843f $X=2.135 $Y=0.805 $X2=0 $Y2=0
cc_267 N_S0_c_231_n N_A3_M1002_g 0.0103041f $X=3.42 $Y=0.18 $X2=0 $Y2=0
cc_268 N_S0_c_231_n N_A1_M1005_g 0.0103041f $X=3.42 $Y=0.18 $X2=0 $Y2=0
cc_269 N_S0_M1001_g N_A1_M1005_g 0.0254677f $X=3.495 $Y=0.805 $X2=0 $Y2=0
cc_270 N_S0_M1011_g N_A1_c_622_n 0.00431314f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_271 N_S0_c_232_n A1 0.0177725f $X=3.495 $Y=1.125 $X2=0 $Y2=0
cc_272 N_S0_c_234_n A1 0.00637639f $X=3.815 $Y=1.46 $X2=0 $Y2=0
cc_273 N_S0_M1011_g A1 0.00294832f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_274 N_S0_c_232_n N_A1_c_624_n 0.0397357f $X=3.495 $Y=1.125 $X2=0 $Y2=0
cc_275 N_S0_c_232_n N_A0_c_673_n 0.00304045f $X=3.495 $Y=1.125 $X2=-0.19
+ $Y2=-0.245
cc_276 N_S0_c_234_n N_A0_c_673_n 0.0539564f $X=3.815 $Y=1.46 $X2=-0.19
+ $Y2=-0.245
cc_277 N_S0_M1011_g N_A0_M1013_g 0.0500919f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_278 N_S0_M1012_g N_VPWR_c_976_n 0.00515681f $X=0.495 $Y=2.74 $X2=0 $Y2=0
cc_279 N_S0_M1011_g N_VPWR_c_978_n 0.001421f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_280 N_S0_M1020_g N_VPWR_c_983_n 0.00390708f $X=1.395 $Y=2.74 $X2=0 $Y2=0
cc_281 N_S0_M1012_g N_VPWR_c_985_n 0.00545712f $X=0.495 $Y=2.74 $X2=0 $Y2=0
cc_282 N_S0_M1011_g N_VPWR_c_986_n 0.00500595f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_283 N_S0_M1012_g N_VPWR_c_975_n 0.00542671f $X=0.495 $Y=2.74 $X2=0 $Y2=0
cc_284 N_S0_M1020_g N_VPWR_c_975_n 0.00542671f $X=1.395 $Y=2.74 $X2=0 $Y2=0
cc_285 N_S0_M1011_g N_VPWR_c_975_n 0.00539454f $X=3.89 $Y=2.73 $X2=0 $Y2=0
cc_286 N_S0_c_242_n N_A_294_506#_c_1073_n 0.00294732f $X=1.395 $Y=2.305 $X2=0
+ $Y2=0
cc_287 N_S0_M1020_g N_A_294_506#_c_1073_n 0.00296302f $X=1.395 $Y=2.74 $X2=0
+ $Y2=0
cc_288 N_S0_c_246_n N_A_294_506#_c_1073_n 0.00621652f $X=1.515 $Y=2.105 $X2=0
+ $Y2=0
cc_289 N_S0_c_242_n N_A_294_506#_c_1065_n 0.00109344f $X=1.395 $Y=2.305 $X2=0
+ $Y2=0
cc_290 N_S0_M1020_g N_A_294_506#_c_1065_n 8.89852e-19 $X=1.395 $Y=2.74 $X2=0
+ $Y2=0
cc_291 N_S0_M1007_g N_A_294_506#_c_1065_n 0.00520728f $X=2.135 $Y=0.805 $X2=0
+ $Y2=0
cc_292 N_S0_c_245_n N_A_294_506#_c_1065_n 0.00546748f $X=1.375 $Y=1.94 $X2=0
+ $Y2=0
cc_293 N_S0_c_246_n N_A_294_506#_c_1065_n 0.0111339f $X=1.515 $Y=2.105 $X2=0
+ $Y2=0
cc_294 S0 N_A_294_506#_c_1065_n 0.00257589f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_295 N_S0_c_231_n N_A_294_506#_c_1068_n 0.00720256f $X=3.42 $Y=0.18 $X2=0
+ $Y2=0
cc_296 N_S0_c_232_n N_A_294_506#_c_1068_n 7.59774e-19 $X=3.495 $Y=1.125 $X2=0
+ $Y2=0
cc_297 N_S0_M1001_g N_A_294_506#_c_1068_n 0.00716554f $X=3.495 $Y=0.805 $X2=0
+ $Y2=0
cc_298 N_S0_c_234_n N_A_294_506#_c_1068_n 0.00333722f $X=3.815 $Y=1.46 $X2=0
+ $Y2=0
cc_299 N_S0_M1007_g N_A_294_506#_c_1069_n 0.00189874f $X=2.135 $Y=0.805 $X2=0
+ $Y2=0
cc_300 N_S0_c_228_n N_A_294_506#_c_1072_n 0.00266209f $X=2.06 $Y=0.18 $X2=0
+ $Y2=0
cc_301 N_S0_M1007_g N_A_294_506#_c_1072_n 0.01154f $X=2.135 $Y=0.805 $X2=0 $Y2=0
cc_302 N_S0_c_231_n N_A_294_506#_c_1072_n 4.626e-19 $X=3.42 $Y=0.18 $X2=0 $Y2=0
cc_303 N_S0_M1011_g N_A_685_504#_c_1196_n 0.00348525f $X=3.89 $Y=2.73 $X2=0
+ $Y2=0
cc_304 N_S0_c_232_n N_A_685_504#_c_1185_n 9.03706e-19 $X=3.495 $Y=1.125 $X2=0
+ $Y2=0
cc_305 N_S0_M1001_g N_A_685_504#_c_1185_n 9.61015e-19 $X=3.495 $Y=0.805 $X2=0
+ $Y2=0
cc_306 N_S0_c_234_n N_A_685_504#_c_1185_n 0.00506474f $X=3.815 $Y=1.46 $X2=0
+ $Y2=0
cc_307 N_S0_M1011_g N_A_685_504#_c_1185_n 4.41403e-19 $X=3.89 $Y=2.73 $X2=0
+ $Y2=0
cc_308 N_S0_M1011_g N_A_685_504#_c_1188_n 0.00616025f $X=3.89 $Y=2.73 $X2=0
+ $Y2=0
cc_309 N_S0_M1011_g N_A_685_504#_c_1189_n 0.00312715f $X=3.89 $Y=2.73 $X2=0
+ $Y2=0
cc_310 N_S0_M1011_g N_A_685_504#_c_1191_n 0.00577222f $X=3.89 $Y=2.73 $X2=0
+ $Y2=0
cc_311 N_S0_M1011_g N_A_685_504#_c_1204_n 0.00590863f $X=3.89 $Y=2.73 $X2=0
+ $Y2=0
cc_312 N_S0_c_232_n N_A_685_504#_c_1205_n 6.79098e-19 $X=3.495 $Y=1.125 $X2=0
+ $Y2=0
cc_313 N_S0_M1001_g N_A_685_504#_c_1205_n 0.00604462f $X=3.495 $Y=0.805 $X2=0
+ $Y2=0
cc_314 N_S0_c_234_n N_A_685_504#_c_1205_n 0.00413524f $X=3.815 $Y=1.46 $X2=0
+ $Y2=0
cc_315 N_S0_M1014_g N_VGND_c_1293_n 0.0251292f $X=0.845 $Y=0.805 $X2=0 $Y2=0
cc_316 N_S0_c_228_n N_VGND_c_1293_n 0.0182681f $X=2.06 $Y=0.18 $X2=0 $Y2=0
cc_317 N_S0_c_229_n N_VGND_c_1293_n 0.00388727f $X=0.92 $Y=0.18 $X2=0 $Y2=0
cc_318 N_S0_M1007_g N_VGND_c_1294_n 0.00608711f $X=2.135 $Y=0.805 $X2=0 $Y2=0
cc_319 N_S0_c_231_n N_VGND_c_1294_n 0.0259687f $X=3.42 $Y=0.18 $X2=0 $Y2=0
cc_320 N_S0_M1001_g N_VGND_c_1294_n 0.00660893f $X=3.495 $Y=0.805 $X2=0 $Y2=0
cc_321 N_S0_c_228_n N_VGND_c_1297_n 0.0463057f $X=2.06 $Y=0.18 $X2=0 $Y2=0
cc_322 N_S0_c_229_n N_VGND_c_1299_n 0.00486043f $X=0.92 $Y=0.18 $X2=0 $Y2=0
cc_323 N_S0_c_231_n N_VGND_c_1300_n 0.0212393f $X=3.42 $Y=0.18 $X2=0 $Y2=0
cc_324 N_S0_c_228_n N_VGND_c_1303_n 0.0329264f $X=2.06 $Y=0.18 $X2=0 $Y2=0
cc_325 N_S0_c_229_n N_VGND_c_1303_n 0.00983503f $X=0.92 $Y=0.18 $X2=0 $Y2=0
cc_326 N_S0_c_231_n N_VGND_c_1303_n 0.047895f $X=3.42 $Y=0.18 $X2=0 $Y2=0
cc_327 N_S0_c_237_n N_VGND_c_1303_n 0.00432083f $X=2.135 $Y=0.18 $X2=0 $Y2=0
cc_328 N_A_31_506#_c_402_n N_A3_M1010_g 0.00689755f $X=2.33 $Y=2.99 $X2=0 $Y2=0
cc_329 N_A_31_506#_c_405_n N_A3_M1010_g 0.00935036f $X=2.415 $Y=2.905 $X2=0
+ $Y2=0
cc_330 N_A_31_506#_c_407_n N_A3_M1010_g 0.00752611f $X=2.5 $Y=2.385 $X2=0 $Y2=0
cc_331 N_A_31_506#_M1009_g N_A3_M1002_g 0.00189267f $X=1.635 $Y=0.805 $X2=0
+ $Y2=0
cc_332 N_A_31_506#_c_395_n N_A3_M1002_g 0.02038f $X=2.055 $Y=1.52 $X2=0 $Y2=0
cc_333 N_A_31_506#_M1004_g A3 2.35688e-19 $X=2.055 $Y=2.73 $X2=0 $Y2=0
cc_334 N_A_31_506#_c_406_n A3 0.0256087f $X=3.275 $Y=2.385 $X2=0 $Y2=0
cc_335 N_A_31_506#_c_407_n A3 0.012371f $X=2.5 $Y=2.385 $X2=0 $Y2=0
cc_336 N_A_31_506#_c_409_n A3 0.00900374f $X=3.535 $Y=2.045 $X2=0 $Y2=0
cc_337 N_A_31_506#_M1004_g N_A3_c_583_n 0.0755527f $X=2.055 $Y=2.73 $X2=0 $Y2=0
cc_338 N_A_31_506#_c_406_n N_A3_c_583_n 0.00443528f $X=3.275 $Y=2.385 $X2=0
+ $Y2=0
cc_339 N_A_31_506#_c_407_n N_A3_c_583_n 2.96179e-19 $X=2.5 $Y=2.385 $X2=0 $Y2=0
cc_340 N_A_31_506#_c_402_n N_A1_M1023_g 3.31545e-19 $X=2.33 $Y=2.99 $X2=0 $Y2=0
cc_341 N_A_31_506#_c_405_n N_A1_M1023_g 0.00107396f $X=2.415 $Y=2.905 $X2=0
+ $Y2=0
cc_342 N_A_31_506#_c_406_n N_A1_M1023_g 0.0138537f $X=3.275 $Y=2.385 $X2=0 $Y2=0
cc_343 N_A_31_506#_c_459_n N_A1_M1023_g 9.28346e-19 $X=3.44 $Y=2.195 $X2=0 $Y2=0
cc_344 N_A_31_506#_c_408_n N_A1_M1023_g 0.0637983f $X=3.44 $Y=2.195 $X2=0 $Y2=0
cc_345 N_A_31_506#_c_409_n N_A1_M1023_g 5.56613e-19 $X=3.535 $Y=2.045 $X2=0
+ $Y2=0
cc_346 N_A_31_506#_c_406_n N_A1_c_622_n 0.00393215f $X=3.275 $Y=2.385 $X2=0
+ $Y2=0
cc_347 N_A_31_506#_c_409_n N_A1_c_622_n 0.00232693f $X=3.535 $Y=2.045 $X2=0
+ $Y2=0
cc_348 N_A_31_506#_c_406_n A1 0.0140129f $X=3.275 $Y=2.385 $X2=0 $Y2=0
cc_349 N_A_31_506#_c_408_n A1 0.00159804f $X=3.44 $Y=2.195 $X2=0 $Y2=0
cc_350 N_A_31_506#_c_409_n A1 0.0236559f $X=3.535 $Y=2.045 $X2=0 $Y2=0
cc_351 N_A_31_506#_c_410_n A1 0.0127335f $X=4.735 $Y=2.075 $X2=0 $Y2=0
cc_352 N_A_31_506#_c_395_n A1 4.51061e-19 $X=2.055 $Y=1.52 $X2=0 $Y2=0
cc_353 N_A_31_506#_c_390_n N_A0_c_673_n 0.0245926f $X=4.83 $Y=1.91 $X2=-0.19
+ $Y2=-0.245
cc_354 N_A_31_506#_c_390_n N_A0_M1013_g 0.00606447f $X=4.83 $Y=1.91 $X2=0 $Y2=0
cc_355 N_A_31_506#_c_410_n N_A0_M1013_g 0.0119731f $X=4.735 $Y=2.075 $X2=0 $Y2=0
cc_356 N_A_31_506#_c_413_n N_A0_M1013_g 0.018402f $X=4.83 $Y=2.075 $X2=0 $Y2=0
cc_357 N_A_31_506#_M1003_g N_A0_c_675_n 0.0416054f $X=3.925 $Y=0.805 $X2=0 $Y2=0
cc_358 N_A_31_506#_c_388_n N_A0_c_675_n 0.0102164f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_359 N_A_31_506#_c_390_n N_A0_c_675_n 0.0128508f $X=4.83 $Y=1.91 $X2=0 $Y2=0
cc_360 N_A_31_506#_c_390_n A0 0.00205617f $X=4.83 $Y=1.91 $X2=0 $Y2=0
cc_361 N_A_31_506#_c_388_n N_A_1029_37#_c_711_n 0.0181329f $X=4.755 $Y=0.18
+ $X2=0 $Y2=0
cc_362 N_A_31_506#_c_390_n N_A_1029_37#_c_715_n 9.96312e-19 $X=4.83 $Y=1.91
+ $X2=0 $Y2=0
cc_363 N_A_31_506#_c_390_n N_A_1029_37#_c_717_n 0.0144023f $X=4.83 $Y=1.91 $X2=0
+ $Y2=0
cc_364 N_A_31_506#_c_410_n N_S1_M1018_g 2.30398e-19 $X=4.735 $Y=2.075 $X2=0
+ $Y2=0
cc_365 N_A_31_506#_c_413_n N_S1_M1018_g 0.0148553f $X=4.83 $Y=2.075 $X2=0 $Y2=0
cc_366 N_A_31_506#_c_390_n N_S1_c_804_n 0.0148553f $X=4.83 $Y=1.91 $X2=0 $Y2=0
cc_367 N_A_31_506#_c_401_n N_VPWR_c_976_n 0.0241757f $X=1.135 $Y=2.445 $X2=0
+ $Y2=0
cc_368 N_A_31_506#_c_403_n N_VPWR_c_976_n 0.0101296f $X=1.305 $Y=2.99 $X2=0
+ $Y2=0
cc_369 N_A_31_506#_M1025_g N_VPWR_c_977_n 0.00149164f $X=3.35 $Y=2.73 $X2=0
+ $Y2=0
cc_370 N_A_31_506#_c_402_n N_VPWR_c_977_n 0.0130135f $X=2.33 $Y=2.99 $X2=0 $Y2=0
cc_371 N_A_31_506#_c_406_n N_VPWR_c_977_n 0.0174569f $X=3.275 $Y=2.385 $X2=0
+ $Y2=0
cc_372 N_A_31_506#_M1004_g N_VPWR_c_983_n 9.59479e-19 $X=2.055 $Y=2.73 $X2=0
+ $Y2=0
cc_373 N_A_31_506#_c_402_n N_VPWR_c_983_n 0.0777206f $X=2.33 $Y=2.99 $X2=0 $Y2=0
cc_374 N_A_31_506#_c_403_n N_VPWR_c_983_n 0.0122334f $X=1.305 $Y=2.99 $X2=0
+ $Y2=0
cc_375 N_A_31_506#_c_400_n N_VPWR_c_985_n 0.00994266f $X=0.28 $Y=2.74 $X2=0
+ $Y2=0
cc_376 N_A_31_506#_M1025_g N_VPWR_c_986_n 0.00563421f $X=3.35 $Y=2.73 $X2=0
+ $Y2=0
cc_377 N_A_31_506#_M1025_g N_VPWR_c_975_n 0.00539454f $X=3.35 $Y=2.73 $X2=0
+ $Y2=0
cc_378 N_A_31_506#_c_400_n N_VPWR_c_975_n 0.0114737f $X=0.28 $Y=2.74 $X2=0 $Y2=0
cc_379 N_A_31_506#_c_401_n N_VPWR_c_975_n 0.0131063f $X=1.135 $Y=2.445 $X2=0
+ $Y2=0
cc_380 N_A_31_506#_c_402_n N_VPWR_c_975_n 0.045054f $X=2.33 $Y=2.99 $X2=0 $Y2=0
cc_381 N_A_31_506#_c_403_n N_VPWR_c_975_n 0.00661802f $X=1.305 $Y=2.99 $X2=0
+ $Y2=0
cc_382 N_A_31_506#_c_406_n N_VPWR_c_975_n 0.0245292f $X=3.275 $Y=2.385 $X2=0
+ $Y2=0
cc_383 N_A_31_506#_c_402_n N_A_294_506#_M1020_d 0.00467726f $X=2.33 $Y=2.99
+ $X2=0 $Y2=0
cc_384 N_A_31_506#_M1004_g N_A_294_506#_c_1073_n 0.0109362f $X=2.055 $Y=2.73
+ $X2=0 $Y2=0
cc_385 N_A_31_506#_c_401_n N_A_294_506#_c_1073_n 0.00372677f $X=1.135 $Y=2.445
+ $X2=0 $Y2=0
cc_386 N_A_31_506#_c_402_n N_A_294_506#_c_1073_n 0.0361387f $X=2.33 $Y=2.99
+ $X2=0 $Y2=0
cc_387 N_A_31_506#_c_405_n N_A_294_506#_c_1073_n 0.00367747f $X=2.415 $Y=2.905
+ $X2=0 $Y2=0
cc_388 N_A_31_506#_M1009_g N_A_294_506#_c_1065_n 0.00205402f $X=1.635 $Y=0.805
+ $X2=0 $Y2=0
cc_389 N_A_31_506#_M1004_g N_A_294_506#_c_1065_n 0.0220394f $X=2.055 $Y=2.73
+ $X2=0 $Y2=0
cc_390 N_A_31_506#_c_393_n N_A_294_506#_c_1065_n 0.0211597f $X=1.485 $Y=1.12
+ $X2=0 $Y2=0
cc_391 N_A_31_506#_c_404_n N_A_294_506#_c_1065_n 0.0218425f $X=1.725 $Y=1.52
+ $X2=0 $Y2=0
cc_392 N_A_31_506#_c_405_n N_A_294_506#_c_1065_n 3.0109e-19 $X=2.415 $Y=2.905
+ $X2=0 $Y2=0
cc_393 N_A_31_506#_c_407_n N_A_294_506#_c_1065_n 0.0143529f $X=2.5 $Y=2.385
+ $X2=0 $Y2=0
cc_394 N_A_31_506#_c_395_n N_A_294_506#_c_1065_n 0.0123485f $X=2.055 $Y=1.52
+ $X2=0 $Y2=0
cc_395 N_A_31_506#_M1003_g N_A_294_506#_c_1068_n 2.47349e-19 $X=3.925 $Y=0.805
+ $X2=0 $Y2=0
cc_396 N_A_31_506#_c_388_n N_A_294_506#_c_1068_n 0.00240993f $X=4.755 $Y=0.18
+ $X2=0 $Y2=0
cc_397 N_A_31_506#_c_390_n N_A_294_506#_c_1068_n 0.0110573f $X=4.83 $Y=1.91
+ $X2=0 $Y2=0
cc_398 N_A_31_506#_M1009_g N_A_294_506#_c_1072_n 0.0070323f $X=1.635 $Y=0.805
+ $X2=0 $Y2=0
cc_399 N_A_31_506#_c_395_n N_A_294_506#_c_1072_n 0.00535124f $X=2.055 $Y=1.52
+ $X2=0 $Y2=0
cc_400 N_A_31_506#_c_402_n A_426_504# 0.00366293f $X=2.33 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_401 N_A_31_506#_M1025_g N_A_685_504#_c_1196_n 0.00236052f $X=3.35 $Y=2.73
+ $X2=0 $Y2=0
cc_402 N_A_31_506#_M1003_g N_A_685_504#_c_1185_n 0.00681803f $X=3.925 $Y=0.805
+ $X2=0 $Y2=0
cc_403 N_A_31_506#_c_410_n N_A_685_504#_c_1188_n 0.0758197f $X=4.735 $Y=2.075
+ $X2=0 $Y2=0
cc_404 N_A_31_506#_c_413_n N_A_685_504#_c_1188_n 0.00892661f $X=4.83 $Y=2.075
+ $X2=0 $Y2=0
cc_405 N_A_31_506#_M1025_g N_A_685_504#_c_1189_n 0.00111961f $X=3.35 $Y=2.73
+ $X2=0 $Y2=0
cc_406 N_A_31_506#_c_406_n N_A_685_504#_c_1189_n 0.0129793f $X=3.275 $Y=2.385
+ $X2=0 $Y2=0
cc_407 N_A_31_506#_c_408_n N_A_685_504#_c_1189_n 2.11399e-19 $X=3.44 $Y=2.195
+ $X2=0 $Y2=0
cc_408 N_A_31_506#_c_410_n N_A_685_504#_c_1189_n 0.0133073f $X=4.735 $Y=2.075
+ $X2=0 $Y2=0
cc_409 N_A_31_506#_c_390_n N_A_685_504#_c_1186_n 0.0129607f $X=4.83 $Y=1.91
+ $X2=0 $Y2=0
cc_410 N_A_31_506#_c_410_n N_A_685_504#_c_1186_n 0.0563899f $X=4.735 $Y=2.075
+ $X2=0 $Y2=0
cc_411 N_A_31_506#_c_413_n N_A_685_504#_c_1186_n 0.00416373f $X=4.83 $Y=2.075
+ $X2=0 $Y2=0
cc_412 N_A_31_506#_c_410_n N_A_685_504#_c_1191_n 0.0121707f $X=4.735 $Y=2.075
+ $X2=0 $Y2=0
cc_413 N_A_31_506#_c_390_n N_A_685_504#_c_1187_n 0.017952f $X=4.83 $Y=1.91 $X2=0
+ $Y2=0
cc_414 N_A_31_506#_c_390_n N_A_685_504#_c_1193_n 0.00661926f $X=4.83 $Y=1.91
+ $X2=0 $Y2=0
cc_415 N_A_31_506#_c_410_n N_A_685_504#_c_1193_n 0.0174453f $X=4.735 $Y=2.075
+ $X2=0 $Y2=0
cc_416 N_A_31_506#_c_406_n N_A_685_504#_c_1204_n 0.00552446f $X=3.275 $Y=2.385
+ $X2=0 $Y2=0
cc_417 N_A_31_506#_c_408_n N_A_685_504#_c_1204_n 0.00199888f $X=3.44 $Y=2.195
+ $X2=0 $Y2=0
cc_418 N_A_31_506#_c_410_n N_A_685_504#_c_1204_n 0.0060962f $X=4.735 $Y=2.075
+ $X2=0 $Y2=0
cc_419 N_A_31_506#_M1003_g N_A_685_504#_c_1205_n 0.00909209f $X=3.925 $Y=0.805
+ $X2=0 $Y2=0
cc_420 N_A_31_506#_M1009_g N_VGND_c_1293_n 0.00153652f $X=1.635 $Y=0.805 $X2=0
+ $Y2=0
cc_421 N_A_31_506#_c_393_n N_VGND_c_1293_n 0.0216087f $X=1.485 $Y=1.12 $X2=0
+ $Y2=0
cc_422 N_A_31_506#_M1003_g N_VGND_c_1295_n 0.00781552f $X=3.925 $Y=0.805 $X2=0
+ $Y2=0
cc_423 N_A_31_506#_c_388_n N_VGND_c_1295_n 0.0248246f $X=4.755 $Y=0.18 $X2=0
+ $Y2=0
cc_424 N_A_31_506#_c_390_n N_VGND_c_1295_n 0.011f $X=4.83 $Y=1.91 $X2=0 $Y2=0
cc_425 N_A_31_506#_c_392_n N_VGND_c_1299_n 0.00466359f $X=0.63 $Y=0.805 $X2=0
+ $Y2=0
cc_426 N_A_31_506#_c_389_n N_VGND_c_1300_n 0.0160075f $X=4 $Y=0.18 $X2=0 $Y2=0
cc_427 N_A_31_506#_c_388_n N_VGND_c_1301_n 0.00932713f $X=4.755 $Y=0.18 $X2=0
+ $Y2=0
cc_428 N_A_31_506#_M1009_g N_VGND_c_1303_n 9.39239e-19 $X=1.635 $Y=0.805 $X2=0
+ $Y2=0
cc_429 N_A_31_506#_c_388_n N_VGND_c_1303_n 0.0309364f $X=4.755 $Y=0.18 $X2=0
+ $Y2=0
cc_430 N_A_31_506#_c_389_n N_VGND_c_1303_n 0.00522251f $X=4 $Y=0.18 $X2=0 $Y2=0
cc_431 N_A_31_506#_c_392_n N_VGND_c_1303_n 0.00760192f $X=0.63 $Y=0.805 $X2=0
+ $Y2=0
cc_432 N_A3_M1010_g N_A1_M1023_g 0.0185464f $X=2.415 $Y=2.73 $X2=0 $Y2=0
cc_433 A3 N_A1_M1023_g 0.00124059f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_434 N_A3_c_583_n N_A1_M1023_g 0.00929883f $X=2.505 $Y=2.035 $X2=0 $Y2=0
cc_435 N_A3_M1002_g N_A1_M1005_g 0.014117f $X=2.495 $Y=0.805 $X2=0 $Y2=0
cc_436 N_A3_M1002_g N_A1_c_622_n 0.00229277f $X=2.495 $Y=0.805 $X2=0 $Y2=0
cc_437 A3 N_A1_c_622_n 0.00105462f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_438 N_A3_c_583_n N_A1_c_622_n 0.00934751f $X=2.505 $Y=2.035 $X2=0 $Y2=0
cc_439 N_A3_M1002_g A1 0.0221489f $X=2.495 $Y=0.805 $X2=0 $Y2=0
cc_440 A3 A1 0.0300257f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_441 N_A3_c_583_n A1 0.00249165f $X=2.505 $Y=2.035 $X2=0 $Y2=0
cc_442 N_A3_M1002_g N_A1_c_624_n 0.0271149f $X=2.495 $Y=0.805 $X2=0 $Y2=0
cc_443 N_A3_M1010_g N_VPWR_c_977_n 0.00159369f $X=2.415 $Y=2.73 $X2=0 $Y2=0
cc_444 N_A3_M1010_g N_VPWR_c_983_n 9.58091e-19 $X=2.415 $Y=2.73 $X2=0 $Y2=0
cc_445 N_A3_M1010_g N_A_294_506#_c_1073_n 3.1532e-19 $X=2.415 $Y=2.73 $X2=0
+ $Y2=0
cc_446 N_A3_M1010_g N_A_294_506#_c_1065_n 5.0079e-19 $X=2.415 $Y=2.73 $X2=0
+ $Y2=0
cc_447 N_A3_M1002_g N_A_294_506#_c_1065_n 0.00738505f $X=2.495 $Y=0.805 $X2=0
+ $Y2=0
cc_448 A3 N_A_294_506#_c_1065_n 0.0147974f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_449 N_A3_c_583_n N_A_294_506#_c_1065_n 0.00521502f $X=2.505 $Y=2.035 $X2=0
+ $Y2=0
cc_450 N_A3_M1002_g N_A_294_506#_c_1068_n 0.0086775f $X=2.495 $Y=0.805 $X2=0
+ $Y2=0
cc_451 N_A3_M1002_g N_A_294_506#_c_1069_n 3.83232e-19 $X=2.495 $Y=0.805 $X2=0
+ $Y2=0
cc_452 N_A3_M1002_g N_A_294_506#_c_1072_n 0.00369786f $X=2.495 $Y=0.805 $X2=0
+ $Y2=0
cc_453 N_A3_M1002_g N_VGND_c_1294_n 0.00864086f $X=2.495 $Y=0.805 $X2=0 $Y2=0
cc_454 N_A3_M1002_g N_VGND_c_1303_n 9.39239e-19 $X=2.495 $Y=0.805 $X2=0 $Y2=0
cc_455 N_A1_M1023_g N_VPWR_c_977_n 0.00830226f $X=2.99 $Y=2.73 $X2=0 $Y2=0
cc_456 N_A1_M1023_g N_VPWR_c_986_n 0.00543288f $X=2.99 $Y=2.73 $X2=0 $Y2=0
cc_457 N_A1_M1023_g N_VPWR_c_975_n 0.00525068f $X=2.99 $Y=2.73 $X2=0 $Y2=0
cc_458 A1 N_A_294_506#_c_1065_n 0.0307984f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_459 N_A1_M1005_g N_A_294_506#_c_1068_n 0.00686339f $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_460 A1 N_A_294_506#_c_1068_n 0.0488832f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_461 A1 N_A_685_504#_c_1185_n 0.0321605f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_462 A1 N_A_685_504#_c_1191_n 0.0145106f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_463 N_A1_M1005_g N_A_685_504#_c_1205_n 0.00103228f $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_464 A1 N_A_685_504#_c_1205_n 0.00855617f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_465 N_A1_M1005_g N_VGND_c_1294_n 0.00973765f $X=3.135 $Y=0.805 $X2=0 $Y2=0
cc_466 A1 N_VGND_c_1294_n 0.0230555f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_467 N_A1_c_624_n N_VGND_c_1294_n 6.95822e-19 $X=3.045 $Y=1.315 $X2=0 $Y2=0
cc_468 N_A1_M1005_g N_VGND_c_1303_n 9.39239e-19 $X=3.135 $Y=0.805 $X2=0 $Y2=0
cc_469 N_A0_M1013_g N_VPWR_c_978_n 0.00986343f $X=4.25 $Y=2.73 $X2=0 $Y2=0
cc_470 N_A0_M1013_g N_VPWR_c_986_n 0.00468165f $X=4.25 $Y=2.73 $X2=0 $Y2=0
cc_471 N_A0_M1013_g N_VPWR_c_975_n 0.00453141f $X=4.25 $Y=2.73 $X2=0 $Y2=0
cc_472 N_A0_c_673_n N_A_294_506#_c_1068_n 0.00536789f $X=4.25 $Y=1.61 $X2=0
+ $Y2=0
cc_473 N_A0_c_675_n N_A_294_506#_c_1068_n 0.00447068f $X=4.285 $Y=1.13 $X2=0
+ $Y2=0
cc_474 A0 N_A_294_506#_c_1068_n 0.0162496f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_475 N_A0_M1013_g N_A_685_504#_c_1196_n 7.60299e-19 $X=4.25 $Y=2.73 $X2=0
+ $Y2=0
cc_476 N_A0_c_673_n N_A_685_504#_c_1185_n 0.00205981f $X=4.25 $Y=1.61 $X2=0
+ $Y2=0
cc_477 N_A0_c_675_n N_A_685_504#_c_1185_n 0.00665536f $X=4.285 $Y=1.13 $X2=0
+ $Y2=0
cc_478 A0 N_A_685_504#_c_1185_n 0.0185483f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_479 N_A0_M1013_g N_A_685_504#_c_1188_n 0.0131775f $X=4.25 $Y=2.73 $X2=0 $Y2=0
cc_480 N_A0_c_673_n N_A_685_504#_c_1186_n 0.00992557f $X=4.25 $Y=1.61 $X2=0
+ $Y2=0
cc_481 N_A0_M1013_g N_A_685_504#_c_1186_n 0.00685186f $X=4.25 $Y=2.73 $X2=0
+ $Y2=0
cc_482 A0 N_A_685_504#_c_1186_n 0.0366657f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_483 N_A0_M1013_g N_A_685_504#_c_1192_n 0.00306478f $X=4.25 $Y=2.73 $X2=0
+ $Y2=0
cc_484 A0 N_A_685_504#_c_1187_n 0.0174674f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_485 N_A0_M1013_g N_A_685_504#_c_1204_n 8.72959e-19 $X=4.25 $Y=2.73 $X2=0
+ $Y2=0
cc_486 N_A0_c_675_n N_A_685_504#_c_1205_n 9.62276e-19 $X=4.285 $Y=1.13 $X2=0
+ $Y2=0
cc_487 N_A0_c_673_n N_VGND_c_1295_n 0.00411873f $X=4.25 $Y=1.61 $X2=0 $Y2=0
cc_488 N_A0_c_675_n N_VGND_c_1295_n 0.00909404f $X=4.285 $Y=1.13 $X2=0 $Y2=0
cc_489 A0 N_VGND_c_1295_n 0.0206119f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_490 N_A0_c_675_n N_VGND_c_1303_n 7.88961e-19 $X=4.285 $Y=1.13 $X2=0 $Y2=0
cc_491 N_A_1029_37#_c_720_n N_S1_M1018_g 0.0326542f $X=5.805 $Y=1.85 $X2=0 $Y2=0
cc_492 N_A_1029_37#_c_713_n N_S1_M1018_g 0.00193246f $X=6.215 $Y=1.69 $X2=0
+ $Y2=0
cc_493 N_A_1029_37#_c_720_n N_S1_c_803_n 0.00611725f $X=5.805 $Y=1.85 $X2=0
+ $Y2=0
cc_494 N_A_1029_37#_c_717_n N_S1_c_804_n 0.010587f $X=5.31 $Y=0.515 $X2=0 $Y2=0
cc_495 N_A_1029_37#_c_711_n N_S1_c_805_n 0.00138059f $X=5.31 $Y=0.35 $X2=0 $Y2=0
cc_496 N_A_1029_37#_c_712_n N_S1_c_805_n 0.00204622f $X=6.4 $Y=1.525 $X2=0 $Y2=0
cc_497 N_A_1029_37#_c_715_n N_S1_c_805_n 0.00595578f $X=6.31 $Y=0.432 $X2=0
+ $Y2=0
cc_498 N_A_1029_37#_c_716_n N_S1_c_805_n 0.002992f $X=6.56 $Y=0.445 $X2=0 $Y2=0
cc_499 N_A_1029_37#_c_717_n N_S1_c_805_n 0.0106755f $X=5.31 $Y=0.515 $X2=0 $Y2=0
cc_500 N_A_1029_37#_c_719_n N_S1_c_806_n 0.00312548f $X=6.05 $Y=1.85 $X2=0 $Y2=0
cc_501 N_A_1029_37#_c_712_n N_S1_c_806_n 0.0133461f $X=6.4 $Y=1.525 $X2=0 $Y2=0
cc_502 N_A_1029_37#_c_713_n N_S1_c_806_n 0.0202106f $X=6.215 $Y=1.69 $X2=0 $Y2=0
cc_503 N_A_1029_37#_c_714_n N_S1_c_806_n 0.00166709f $X=6.4 $Y=1.69 $X2=0 $Y2=0
cc_504 N_A_1029_37#_c_715_n N_S1_c_806_n 0.00429467f $X=6.31 $Y=0.432 $X2=0
+ $Y2=0
cc_505 N_A_1029_37#_c_716_n N_S1_c_806_n 0.00396731f $X=6.56 $Y=0.445 $X2=0
+ $Y2=0
cc_506 N_A_1029_37#_c_713_n N_S1_M1022_g 0.00539025f $X=6.215 $Y=1.69 $X2=0
+ $Y2=0
cc_507 N_A_1029_37#_c_714_n N_S1_M1022_g 7.25655e-19 $X=6.4 $Y=1.69 $X2=0 $Y2=0
cc_508 N_A_1029_37#_c_723_n N_S1_M1022_g 0.00479831f $X=6.465 $Y=2.225 $X2=0
+ $Y2=0
cc_509 N_A_1029_37#_c_724_n N_S1_M1022_g 0.00501741f $X=6.465 $Y=2.06 $X2=0
+ $Y2=0
cc_510 N_A_1029_37#_c_712_n N_S1_M1021_g 0.00753272f $X=6.4 $Y=1.525 $X2=0 $Y2=0
cc_511 N_A_1029_37#_c_719_n N_S1_c_808_n 0.00611725f $X=6.05 $Y=1.85 $X2=0 $Y2=0
cc_512 N_A_1029_37#_c_712_n N_S1_c_808_n 0.00149528f $X=6.4 $Y=1.525 $X2=0 $Y2=0
cc_513 N_A_1029_37#_c_713_n N_S1_c_808_n 0.00209298f $X=6.215 $Y=1.69 $X2=0
+ $Y2=0
cc_514 N_A_1029_37#_c_715_n N_S1_c_808_n 6.0795e-19 $X=6.31 $Y=0.432 $X2=0 $Y2=0
cc_515 N_A_1029_37#_c_717_n N_S1_c_808_n 9.02921e-19 $X=5.31 $Y=0.515 $X2=0
+ $Y2=0
cc_516 N_A_1029_37#_c_712_n S1 0.0579754f $X=6.4 $Y=1.525 $X2=0 $Y2=0
cc_517 N_A_1029_37#_c_713_n S1 2.67214e-19 $X=6.215 $Y=1.69 $X2=0 $Y2=0
cc_518 N_A_1029_37#_c_714_n S1 0.0245222f $X=6.4 $Y=1.69 $X2=0 $Y2=0
cc_519 N_A_1029_37#_c_712_n N_S1_c_811_n 0.00534349f $X=6.4 $Y=1.525 $X2=0 $Y2=0
cc_520 N_A_1029_37#_c_713_n N_S1_c_811_n 0.0185793f $X=6.215 $Y=1.69 $X2=0 $Y2=0
cc_521 N_A_1029_37#_c_714_n N_S1_c_811_n 0.00196112f $X=6.4 $Y=1.69 $X2=0 $Y2=0
cc_522 N_A_1029_37#_c_720_n N_A_1075_493#_c_903_n 0.00604102f $X=5.805 $Y=1.85
+ $X2=0 $Y2=0
cc_523 N_A_1029_37#_c_711_n N_A_1075_493#_c_914_n 0.00115213f $X=5.31 $Y=0.35
+ $X2=0 $Y2=0
cc_524 N_A_1029_37#_c_715_n N_A_1075_493#_c_914_n 0.0142221f $X=6.31 $Y=0.432
+ $X2=0 $Y2=0
cc_525 N_A_1029_37#_c_717_n N_A_1075_493#_c_914_n 0.00124796f $X=5.31 $Y=0.515
+ $X2=0 $Y2=0
cc_526 N_A_1029_37#_M1000_g N_A_1075_493#_c_910_n 4.95435e-19 $X=5.73 $Y=2.675
+ $X2=0 $Y2=0
cc_527 N_A_1029_37#_c_723_n N_A_1075_493#_c_910_n 0.00752331f $X=6.465 $Y=2.225
+ $X2=0 $Y2=0
cc_528 N_A_1029_37#_M1000_g N_A_1075_493#_c_911_n 0.01286f $X=5.73 $Y=2.675
+ $X2=0 $Y2=0
cc_529 N_A_1029_37#_c_723_n N_A_1075_493#_c_911_n 0.00421457f $X=6.465 $Y=2.225
+ $X2=0 $Y2=0
cc_530 N_A_1029_37#_M1000_g N_A_1075_493#_c_912_n 0.00292875f $X=5.73 $Y=2.675
+ $X2=0 $Y2=0
cc_531 N_A_1029_37#_c_723_n N_A_1075_493#_c_912_n 0.00362047f $X=6.465 $Y=2.225
+ $X2=0 $Y2=0
cc_532 N_A_1029_37#_M1000_g N_VPWR_c_979_n 8.16603e-19 $X=5.73 $Y=2.675 $X2=0
+ $Y2=0
cc_533 N_A_1029_37#_c_724_n N_VPWR_c_981_n 0.00205926f $X=6.465 $Y=2.06 $X2=0
+ $Y2=0
cc_534 N_A_1029_37#_c_719_n N_A_294_506#_c_1066_n 0.0021367f $X=6.05 $Y=1.85
+ $X2=0 $Y2=0
cc_535 N_A_1029_37#_c_713_n N_A_294_506#_c_1066_n 0.00200338f $X=6.215 $Y=1.69
+ $X2=0 $Y2=0
cc_536 N_A_1029_37#_c_714_n N_A_294_506#_c_1066_n 0.00147574f $X=6.4 $Y=1.69
+ $X2=0 $Y2=0
cc_537 N_A_1029_37#_c_715_n N_A_294_506#_c_1066_n 2.72334e-19 $X=6.31 $Y=0.432
+ $X2=0 $Y2=0
cc_538 N_A_1029_37#_M1000_g N_A_294_506#_c_1075_n 0.00310761f $X=5.73 $Y=2.675
+ $X2=0 $Y2=0
cc_539 N_A_1029_37#_c_719_n N_A_294_506#_c_1075_n 0.00410483f $X=6.05 $Y=1.85
+ $X2=0 $Y2=0
cc_540 N_A_1029_37#_M1000_g N_A_294_506#_c_1067_n 0.0149575f $X=5.73 $Y=2.675
+ $X2=0 $Y2=0
cc_541 N_A_1029_37#_c_719_n N_A_294_506#_c_1067_n 0.0107784f $X=6.05 $Y=1.85
+ $X2=0 $Y2=0
cc_542 N_A_1029_37#_c_720_n N_A_294_506#_c_1067_n 0.00175013f $X=5.805 $Y=1.85
+ $X2=0 $Y2=0
cc_543 N_A_1029_37#_c_712_n N_A_294_506#_c_1067_n 0.00585216f $X=6.4 $Y=1.525
+ $X2=0 $Y2=0
cc_544 N_A_1029_37#_c_713_n N_A_294_506#_c_1067_n 0.00279606f $X=6.215 $Y=1.69
+ $X2=0 $Y2=0
cc_545 N_A_1029_37#_c_714_n N_A_294_506#_c_1067_n 0.0246931f $X=6.4 $Y=1.69
+ $X2=0 $Y2=0
cc_546 N_A_1029_37#_c_724_n N_A_294_506#_c_1067_n 0.0247573f $X=6.465 $Y=2.06
+ $X2=0 $Y2=0
cc_547 N_A_1029_37#_c_711_n N_A_294_506#_c_1068_n 4.23553e-19 $X=5.31 $Y=0.35
+ $X2=0 $Y2=0
cc_548 N_A_1029_37#_c_715_n N_A_294_506#_c_1068_n 0.0127369f $X=6.31 $Y=0.432
+ $X2=0 $Y2=0
cc_549 N_A_1029_37#_c_717_n N_A_294_506#_c_1068_n 0.00412651f $X=5.31 $Y=0.515
+ $X2=0 $Y2=0
cc_550 N_A_1029_37#_c_712_n N_A_294_506#_c_1070_n 0.00727882f $X=6.4 $Y=1.525
+ $X2=0 $Y2=0
cc_551 N_A_1029_37#_c_714_n N_A_294_506#_c_1070_n 2.76875e-19 $X=6.4 $Y=1.69
+ $X2=0 $Y2=0
cc_552 N_A_1029_37#_c_715_n N_A_294_506#_c_1070_n 0.00183845f $X=6.31 $Y=0.432
+ $X2=0 $Y2=0
cc_553 N_A_1029_37#_c_712_n N_A_294_506#_c_1071_n 0.0496418f $X=6.4 $Y=1.525
+ $X2=0 $Y2=0
cc_554 N_A_1029_37#_c_715_n N_A_294_506#_c_1071_n 0.0223373f $X=6.31 $Y=0.432
+ $X2=0 $Y2=0
cc_555 N_A_1029_37#_c_711_n N_A_685_504#_c_1187_n 0.00230673f $X=5.31 $Y=0.35
+ $X2=0 $Y2=0
cc_556 N_A_1029_37#_c_715_n N_A_685_504#_c_1187_n 0.00547799f $X=6.31 $Y=0.432
+ $X2=0 $Y2=0
cc_557 N_A_1029_37#_c_717_n N_A_685_504#_c_1187_n 0.00148021f $X=5.31 $Y=0.515
+ $X2=0 $Y2=0
cc_558 N_A_1029_37#_c_711_n N_VGND_c_1295_n 8.45456e-19 $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_559 N_A_1029_37#_c_715_n N_VGND_c_1295_n 0.00929837f $X=6.31 $Y=0.432 $X2=0
+ $Y2=0
cc_560 N_A_1029_37#_c_711_n N_VGND_c_1301_n 0.00647615f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_561 N_A_1029_37#_c_715_n N_VGND_c_1301_n 0.0999503f $X=6.31 $Y=0.432 $X2=0
+ $Y2=0
cc_562 N_A_1029_37#_M1021_s N_VGND_c_1303_n 0.00221698f $X=6.435 $Y=0.235 $X2=0
+ $Y2=0
cc_563 N_A_1029_37#_c_711_n N_VGND_c_1303_n 0.00945174f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_564 N_A_1029_37#_c_715_n N_VGND_c_1303_n 0.0571676f $X=6.31 $Y=0.432 $X2=0
+ $Y2=0
cc_565 N_S1_M1021_g N_A_1075_493#_c_900_n 0.018639f $X=6.775 $Y=0.445 $X2=0
+ $Y2=0
cc_566 S1 N_A_1075_493#_c_901_n 0.0011565f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_567 N_S1_M1021_g N_A_1075_493#_c_902_n 0.00831755f $X=6.775 $Y=0.445 $X2=0
+ $Y2=0
cc_568 N_S1_c_809_n N_A_1075_493#_c_902_n 0.0294617f $X=6.755 $Y=1.23 $X2=0
+ $Y2=0
cc_569 S1 N_A_1075_493#_c_902_n 0.00635654f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_570 N_S1_M1022_g N_A_1075_493#_c_907_n 0.0113077f $X=6.68 $Y=2.225 $X2=0
+ $Y2=0
cc_571 N_S1_c_814_n N_A_1075_493#_c_907_n 0.00413581f $X=6.755 $Y=1.825 $X2=0
+ $Y2=0
cc_572 S1 N_A_1075_493#_c_907_n 5.24125e-19 $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_573 N_S1_M1018_g N_A_1075_493#_c_903_n 0.00821168f $X=5.3 $Y=2.675 $X2=0
+ $Y2=0
cc_574 N_S1_c_803_n N_A_1075_493#_c_903_n 0.0156376f $X=5.66 $Y=1.49 $X2=0 $Y2=0
cc_575 N_S1_c_805_n N_A_1075_493#_c_903_n 9.73062e-19 $X=5.76 $Y=1.155 $X2=0
+ $Y2=0
cc_576 N_S1_c_808_n N_A_1075_493#_c_903_n 0.00657009f $X=5.747 $Y=1.23 $X2=0
+ $Y2=0
cc_577 N_S1_M1018_g N_A_1075_493#_c_909_n 0.00352394f $X=5.3 $Y=2.675 $X2=0
+ $Y2=0
cc_578 N_S1_c_803_n N_A_1075_493#_c_914_n 6.64275e-19 $X=5.66 $Y=1.49 $X2=0
+ $Y2=0
cc_579 N_S1_M1022_g N_A_1075_493#_c_910_n 9.99569e-19 $X=6.68 $Y=2.225 $X2=0
+ $Y2=0
cc_580 N_S1_M1022_g N_A_1075_493#_c_912_n 0.0103162f $X=6.68 $Y=2.225 $X2=0
+ $Y2=0
cc_581 N_S1_M1018_g N_VPWR_c_978_n 0.0038491f $X=5.3 $Y=2.675 $X2=0 $Y2=0
cc_582 N_S1_M1018_g N_VPWR_c_979_n 0.00502202f $X=5.3 $Y=2.675 $X2=0 $Y2=0
cc_583 N_S1_M1022_g N_VPWR_c_980_n 0.0027316f $X=6.68 $Y=2.225 $X2=0 $Y2=0
cc_584 N_S1_M1022_g N_VPWR_c_981_n 0.00153902f $X=6.68 $Y=2.225 $X2=0 $Y2=0
cc_585 N_S1_c_814_n N_VPWR_c_981_n 9.21813e-19 $X=6.755 $Y=1.825 $X2=0 $Y2=0
cc_586 S1 N_VPWR_c_981_n 0.0268617f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_587 N_S1_M1018_g N_VPWR_c_975_n 0.0052212f $X=5.3 $Y=2.675 $X2=0 $Y2=0
cc_588 N_S1_c_806_n N_A_294_506#_c_1066_n 0.00744524f $X=6.59 $Y=1.23 $X2=0
+ $Y2=0
cc_589 N_S1_c_808_n N_A_294_506#_c_1066_n 0.00380138f $X=5.747 $Y=1.23 $X2=0
+ $Y2=0
cc_590 N_S1_M1022_g N_A_294_506#_c_1075_n 0.00276976f $X=6.68 $Y=2.225 $X2=0
+ $Y2=0
cc_591 N_S1_c_808_n N_A_294_506#_c_1067_n 0.00714154f $X=5.747 $Y=1.23 $X2=0
+ $Y2=0
cc_592 N_S1_c_811_n N_A_294_506#_c_1067_n 2.47116e-19 $X=6.755 $Y=1.32 $X2=0
+ $Y2=0
cc_593 N_S1_c_803_n N_A_294_506#_c_1068_n 6.3154e-19 $X=5.66 $Y=1.49 $X2=0 $Y2=0
cc_594 N_S1_c_804_n N_A_294_506#_c_1068_n 8.29737e-19 $X=5.375 $Y=1.49 $X2=0
+ $Y2=0
cc_595 N_S1_c_805_n N_A_294_506#_c_1068_n 0.00541524f $X=5.76 $Y=1.155 $X2=0
+ $Y2=0
cc_596 N_S1_c_808_n N_A_294_506#_c_1068_n 6.20255e-19 $X=5.747 $Y=1.23 $X2=0
+ $Y2=0
cc_597 N_S1_c_805_n N_A_294_506#_c_1071_n 0.0073876f $X=5.76 $Y=1.155 $X2=0
+ $Y2=0
cc_598 N_S1_c_806_n N_A_294_506#_c_1071_n 0.00560041f $X=6.59 $Y=1.23 $X2=0
+ $Y2=0
cc_599 N_S1_c_808_n N_A_294_506#_c_1071_n 2.17867e-19 $X=5.747 $Y=1.23 $X2=0
+ $Y2=0
cc_600 N_S1_M1018_g N_A_685_504#_c_1192_n 0.00376335f $X=5.3 $Y=2.675 $X2=0
+ $Y2=0
cc_601 N_S1_c_804_n N_A_685_504#_c_1187_n 0.00451592f $X=5.375 $Y=1.49 $X2=0
+ $Y2=0
cc_602 N_S1_M1018_g N_A_685_504#_c_1193_n 0.0123884f $X=5.3 $Y=2.675 $X2=0 $Y2=0
cc_603 N_S1_M1018_g N_A_685_504#_c_1194_n 0.0053532f $X=5.3 $Y=2.675 $X2=0 $Y2=0
cc_604 N_S1_M1018_g N_A_685_504#_c_1195_n 0.00390261f $X=5.3 $Y=2.675 $X2=0
+ $Y2=0
cc_605 N_S1_M1022_g N_X_c_1275_n 3.53152e-19 $X=6.68 $Y=2.225 $X2=0 $Y2=0
cc_606 N_S1_M1021_g N_X_c_1275_n 3.33905e-19 $X=6.775 $Y=0.445 $X2=0 $Y2=0
cc_607 N_S1_c_809_n N_X_c_1275_n 4.95397e-19 $X=6.755 $Y=1.23 $X2=0 $Y2=0
cc_608 S1 N_X_c_1275_n 0.0842087f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_609 N_S1_M1021_g N_VGND_c_1296_n 0.00315529f $X=6.775 $Y=0.445 $X2=0 $Y2=0
cc_610 S1 N_VGND_c_1296_n 0.0186433f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_611 N_S1_c_805_n N_VGND_c_1301_n 5.34712e-19 $X=5.76 $Y=1.155 $X2=0 $Y2=0
cc_612 N_S1_M1021_g N_VGND_c_1301_n 0.00585385f $X=6.775 $Y=0.445 $X2=0 $Y2=0
cc_613 N_S1_M1021_g N_VGND_c_1303_n 0.00756476f $X=6.775 $Y=0.445 $X2=0 $Y2=0
cc_614 S1 N_VGND_c_1303_n 0.00696804f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_615 N_A_1075_493#_c_904_n N_VPWR_c_979_n 0.00344245f $X=7.13 $Y=2.855 $X2=0
+ $Y2=0
cc_616 N_A_1075_493#_c_909_n N_VPWR_c_979_n 0.0135481f $X=5.61 $Y=2.99 $X2=0
+ $Y2=0
cc_617 N_A_1075_493#_c_911_n N_VPWR_c_979_n 0.0728606f $X=6.415 $Y=2.927 $X2=0
+ $Y2=0
cc_618 N_A_1075_493#_c_912_n N_VPWR_c_979_n 0.00582945f $X=6.58 $Y=2.855 $X2=0
+ $Y2=0
cc_619 N_A_1075_493#_c_904_n N_VPWR_c_980_n 0.00307725f $X=7.13 $Y=2.855 $X2=0
+ $Y2=0
cc_620 N_A_1075_493#_M1019_g N_VPWR_c_980_n 4.5639e-19 $X=7.205 $Y=2.335 $X2=0
+ $Y2=0
cc_621 N_A_1075_493#_M1019_g N_VPWR_c_981_n 0.00187421f $X=7.205 $Y=2.335 $X2=0
+ $Y2=0
cc_622 N_A_1075_493#_c_904_n N_VPWR_c_982_n 0.0185011f $X=7.13 $Y=2.855 $X2=0
+ $Y2=0
cc_623 N_A_1075_493#_M1019_g N_VPWR_c_982_n 0.00415414f $X=7.205 $Y=2.335 $X2=0
+ $Y2=0
cc_624 N_A_1075_493#_c_910_n N_VPWR_c_982_n 0.0224062f $X=6.58 $Y=2.945 $X2=0
+ $Y2=0
cc_625 N_A_1075_493#_c_912_n N_VPWR_c_982_n 0.00214924f $X=6.58 $Y=2.855 $X2=0
+ $Y2=0
cc_626 N_A_1075_493#_c_904_n N_VPWR_c_987_n 0.00554211f $X=7.13 $Y=2.855 $X2=0
+ $Y2=0
cc_627 N_A_1075_493#_c_904_n N_VPWR_c_975_n 0.0104015f $X=7.13 $Y=2.855 $X2=0
+ $Y2=0
cc_628 N_A_1075_493#_c_909_n N_VPWR_c_975_n 0.0073762f $X=5.61 $Y=2.99 $X2=0
+ $Y2=0
cc_629 N_A_1075_493#_c_911_n N_VPWR_c_975_n 0.0413111f $X=6.415 $Y=2.927 $X2=0
+ $Y2=0
cc_630 N_A_1075_493#_c_912_n N_VPWR_c_975_n 0.00834335f $X=6.58 $Y=2.855 $X2=0
+ $Y2=0
cc_631 N_A_1075_493#_c_903_n N_A_294_506#_c_1066_n 0.104807f $X=5.515 $Y=2.74
+ $X2=0 $Y2=0
cc_632 N_A_1075_493#_c_911_n N_A_294_506#_c_1075_n 0.0222155f $X=6.415 $Y=2.927
+ $X2=0 $Y2=0
cc_633 N_A_1075_493#_M1016_d N_A_294_506#_c_1068_n 0.0014777f $X=5.405 $Y=0.625
+ $X2=0 $Y2=0
cc_634 N_A_1075_493#_c_914_n N_A_294_506#_c_1068_n 0.0152016f $X=5.545 $Y=0.835
+ $X2=0 $Y2=0
cc_635 N_A_1075_493#_c_903_n N_A_294_506#_c_1070_n 2.30567e-19 $X=5.515 $Y=2.74
+ $X2=0 $Y2=0
cc_636 N_A_1075_493#_c_914_n N_A_294_506#_c_1070_n 3.75261e-19 $X=5.545 $Y=0.835
+ $X2=0 $Y2=0
cc_637 N_A_1075_493#_c_903_n N_A_294_506#_c_1071_n 0.0110152f $X=5.515 $Y=2.74
+ $X2=0 $Y2=0
cc_638 N_A_1075_493#_c_914_n N_A_294_506#_c_1071_n 0.0143737f $X=5.545 $Y=0.835
+ $X2=0 $Y2=0
cc_639 N_A_1075_493#_c_914_n N_A_685_504#_c_1187_n 0.0445917f $X=5.545 $Y=0.835
+ $X2=0 $Y2=0
cc_640 N_A_1075_493#_c_903_n N_A_685_504#_c_1193_n 0.0440129f $X=5.515 $Y=2.74
+ $X2=0 $Y2=0
cc_641 N_A_1075_493#_c_903_n N_A_685_504#_c_1194_n 0.0123101f $X=5.515 $Y=2.74
+ $X2=0 $Y2=0
cc_642 N_A_1075_493#_c_903_n N_A_685_504#_c_1195_n 0.0136324f $X=5.515 $Y=2.74
+ $X2=0 $Y2=0
cc_643 N_A_1075_493#_M1019_g N_X_c_1275_n 0.00488989f $X=7.205 $Y=2.335 $X2=0
+ $Y2=0
cc_644 N_A_1075_493#_c_900_n N_X_c_1275_n 0.00509062f $X=7.22 $Y=0.765 $X2=0
+ $Y2=0
cc_645 N_A_1075_493#_c_901_n N_X_c_1275_n 0.00525309f $X=7.22 $Y=0.915 $X2=0
+ $Y2=0
cc_646 N_A_1075_493#_c_902_n N_X_c_1275_n 0.0250333f $X=7.22 $Y=1.755 $X2=0
+ $Y2=0
cc_647 N_A_1075_493#_c_907_n N_X_c_1275_n 0.00593199f $X=7.22 $Y=1.905 $X2=0
+ $Y2=0
cc_648 N_A_1075_493#_c_900_n N_VGND_c_1296_n 0.0031247f $X=7.22 $Y=0.765 $X2=0
+ $Y2=0
cc_649 N_A_1075_493#_c_900_n N_VGND_c_1302_n 0.00585385f $X=7.22 $Y=0.765 $X2=0
+ $Y2=0
cc_650 N_A_1075_493#_c_900_n N_VGND_c_1303_n 0.0117828f $X=7.22 $Y=0.765 $X2=0
+ $Y2=0
cc_651 N_VPWR_c_978_n N_A_685_504#_c_1188_n 0.0238095f $X=4.465 $Y=2.775 $X2=0
+ $Y2=0
cc_652 N_VPWR_c_975_n N_A_685_504#_c_1188_n 0.0252952f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_653 N_VPWR_c_978_n N_A_685_504#_c_1192_n 0.00977198f $X=4.465 $Y=2.775 $X2=0
+ $Y2=0
cc_654 N_VPWR_c_979_n N_A_685_504#_c_1192_n 0.00815216f $X=6.915 $Y=3.33 $X2=0
+ $Y2=0
cc_655 N_VPWR_c_975_n N_A_685_504#_c_1192_n 0.0109491f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_978_n N_A_685_504#_c_1204_n 0.00910001f $X=4.465 $Y=2.775 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_986_n N_A_685_504#_c_1204_n 0.0124424f $X=4.3 $Y=3.33 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_975_n N_A_685_504#_c_1204_n 0.0143991f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_980_n N_X_c_1275_n 0.00141149f $X=6.947 $Y=2.468 $X2=0 $Y2=0
cc_660 N_VPWR_c_981_n N_X_c_1275_n 0.00143894f $X=6.895 $Y=2.16 $X2=0 $Y2=0
cc_661 N_VPWR_c_987_n N_X_c_1275_n 0.00579333f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_662 N_VPWR_c_975_n N_X_c_1275_n 0.00891079f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_663 N_A_294_506#_c_1068_n N_A_685_504#_M1001_d 0.00363728f $X=5.855 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_664 N_A_294_506#_c_1068_n N_A_685_504#_c_1185_n 0.00839562f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_665 N_A_294_506#_c_1068_n N_A_685_504#_c_1186_n 0.0121509f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_666 N_A_294_506#_c_1068_n N_A_685_504#_c_1187_n 0.034262f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_667 N_A_294_506#_c_1068_n N_A_685_504#_c_1205_n 0.0362318f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_668 N_A_294_506#_c_1068_n N_VGND_M1002_d 0.00672387f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_669 N_A_294_506#_c_1068_n N_VGND_M1024_d 0.00203297f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_670 N_A_294_506#_c_1072_n N_VGND_c_1293_n 0.0066936f $X=2.075 $Y=0.827 $X2=0
+ $Y2=0
cc_671 N_A_294_506#_c_1068_n N_VGND_c_1294_n 0.019146f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_672 N_A_294_506#_c_1069_n N_VGND_c_1294_n 3.24904e-19 $X=2.305 $Y=0.925 $X2=0
+ $Y2=0
cc_673 N_A_294_506#_c_1072_n N_VGND_c_1294_n 0.014582f $X=2.075 $Y=0.827 $X2=0
+ $Y2=0
cc_674 N_A_294_506#_c_1068_n N_VGND_c_1295_n 0.0180367f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_675 N_A_294_506#_c_1072_n N_VGND_c_1297_n 0.00801408f $X=2.075 $Y=0.827 $X2=0
+ $Y2=0
cc_676 N_A_294_506#_c_1072_n N_VGND_c_1303_n 0.0126297f $X=2.075 $Y=0.827 $X2=0
+ $Y2=0
cc_677 N_A_294_506#_c_1068_n A_442_119# 0.00533292f $X=5.855 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_678 N_A_294_506#_c_1072_n A_442_119# 0.00647728f $X=2.075 $Y=0.827 $X2=-0.19
+ $Y2=-0.245
cc_679 N_A_294_506#_c_1068_n A_642_119# 0.0072202f $X=5.855 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_680 N_A_294_506#_c_1068_n A_800_119# 0.00642416f $X=5.855 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_681 N_A_685_504#_c_1205_n N_VGND_c_1294_n 0.00837955f $X=3.95 $Y=0.805 $X2=0
+ $Y2=0
cc_682 N_A_685_504#_c_1187_n N_VGND_c_1295_n 0.0156405f $X=5.115 $Y=0.835 $X2=0
+ $Y2=0
cc_683 N_A_685_504#_c_1205_n N_VGND_c_1295_n 0.00824646f $X=3.95 $Y=0.805 $X2=0
+ $Y2=0
cc_684 N_A_685_504#_c_1205_n N_VGND_c_1300_n 0.00737045f $X=3.95 $Y=0.805 $X2=0
+ $Y2=0
cc_685 N_A_685_504#_c_1187_n N_VGND_c_1301_n 0.0035101f $X=5.115 $Y=0.835 $X2=0
+ $Y2=0
cc_686 N_A_685_504#_c_1187_n N_VGND_c_1303_n 0.00598891f $X=5.115 $Y=0.835 $X2=0
+ $Y2=0
cc_687 N_A_685_504#_c_1205_n N_VGND_c_1303_n 0.0132602f $X=3.95 $Y=0.805 $X2=0
+ $Y2=0
cc_688 N_X_c_1275_n N_VGND_c_1302_n 0.0165868f $X=7.42 $Y=0.445 $X2=0 $Y2=0
cc_689 N_X_M1008_d N_VGND_c_1303_n 0.00223914f $X=7.28 $Y=0.235 $X2=0 $Y2=0
cc_690 N_X_c_1275_n N_VGND_c_1303_n 0.0114448f $X=7.42 $Y=0.445 $X2=0 $Y2=0
