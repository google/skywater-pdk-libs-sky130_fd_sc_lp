* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buflp_m A VGND VNB VPB VPWR X
X0 a_120_120# a_90_94# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_90_94# a_120_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_304_490# A a_90_94# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR A a_304_490# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 X a_90_94# a_120_490# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND A a_278_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_120_490# a_90_94# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_278_120# A a_90_94# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
