* File: sky130_fd_sc_lp__xor2_0.pxi.spice
* Created: Fri Aug 28 11:36:04 2020
* 
x_PM_SKY130_FD_SC_LP__XOR2_0%B N_B_M1001_g N_B_M1009_g N_B_M1006_g N_B_M1005_g
+ N_B_c_74_n N_B_c_75_n N_B_c_76_n B B B B N_B_c_78_n N_B_c_79_n
+ PM_SKY130_FD_SC_LP__XOR2_0%B
x_PM_SKY130_FD_SC_LP__XOR2_0%A N_A_M1003_g N_A_M1002_g N_A_M1000_g N_A_M1004_g
+ N_A_c_156_n N_A_c_151_n A A N_A_c_153_n PM_SKY130_FD_SC_LP__XOR2_0%A
x_PM_SKY130_FD_SC_LP__XOR2_0%A_27_481# N_A_27_481#_M1009_d N_A_27_481#_M1001_s
+ N_A_27_481#_c_201_n N_A_27_481#_c_202_n N_A_27_481#_c_203_n
+ N_A_27_481#_M1008_g N_A_27_481#_M1007_g N_A_27_481#_c_205_n
+ N_A_27_481#_c_214_n N_A_27_481#_c_215_n N_A_27_481#_c_216_n
+ N_A_27_481#_c_206_n N_A_27_481#_c_207_n N_A_27_481#_c_208_n
+ N_A_27_481#_c_209_n N_A_27_481#_c_210_n N_A_27_481#_c_211_n
+ N_A_27_481#_c_212_n PM_SKY130_FD_SC_LP__XOR2_0%A_27_481#
x_PM_SKY130_FD_SC_LP__XOR2_0%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_c_285_n
+ N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n
+ VPWR N_VPWR_c_291_n N_VPWR_c_284_n PM_SKY130_FD_SC_LP__XOR2_0%VPWR
x_PM_SKY130_FD_SC_LP__XOR2_0%A_274_481# N_A_274_481#_M1000_d
+ N_A_274_481#_M1007_d N_A_274_481#_c_323_n N_A_274_481#_c_324_n
+ N_A_274_481#_c_325_n N_A_274_481#_c_326_n N_A_274_481#_c_327_n
+ N_A_274_481#_c_328_n PM_SKY130_FD_SC_LP__XOR2_0%A_274_481#
x_PM_SKY130_FD_SC_LP__XOR2_0%X N_X_M1005_d N_X_M1007_s N_X_c_357_n N_X_c_358_n
+ N_X_c_354_n N_X_c_355_n X X N_X_c_356_n X PM_SKY130_FD_SC_LP__XOR2_0%X
x_PM_SKY130_FD_SC_LP__XOR2_0%VGND N_VGND_M1009_s N_VGND_M1002_d N_VGND_M1008_d
+ N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n
+ N_VGND_c_392_n VGND N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n
+ PM_SKY130_FD_SC_LP__XOR2_0%VGND
cc_1 VNB N_B_M1009_g 0.039103f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.635
cc_2 VNB N_B_M1005_g 0.0482842f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.635
cc_3 VNB N_B_c_74_n 0.00366547f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.565
cc_4 VNB N_B_c_75_n 0.00504029f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.35
cc_5 VNB N_B_c_76_n 0.0675301f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.35
cc_6 VNB B 0.00493211f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_7 VNB N_B_c_78_n 0.0155732f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.685
cc_8 VNB N_B_c_79_n 0.00422266f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.71
cc_9 VNB N_A_M1002_g 0.0235133f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.635
cc_10 VNB N_A_M1004_g 0.0228421f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.635
cc_11 VNB N_A_c_151_n 0.0226249f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_12 VNB A 0.00527543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_c_153_n 0.0283751f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.35
cc_14 VNB N_A_27_481#_c_201_n 0.0134481f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.635
cc_15 VNB N_A_27_481#_c_202_n 0.0163206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_481#_c_203_n 0.0246214f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=1.85
cc_17 VNB N_A_27_481#_M1007_g 0.0417824f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.635
cc_18 VNB N_A_27_481#_c_205_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.565
cc_19 VNB N_A_27_481#_c_206_n 0.00319953f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB N_A_27_481#_c_207_n 0.0302706f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_21 VNB N_A_27_481#_c_208_n 0.00452216f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_22 VNB N_A_27_481#_c_209_n 0.00380992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_481#_c_210_n 0.043839f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.35
cc_24 VNB N_A_27_481#_c_211_n 4.41111e-19 $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.69
cc_25 VNB N_A_27_481#_c_212_n 0.00500661f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.855
cc_26 VNB N_VPWR_c_284_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.185
cc_27 VNB N_X_c_354_n 0.00147068f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.725
cc_28 VNB N_X_c_355_n 0.00433043f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.52
cc_29 VNB N_X_c_356_n 0.00649516f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.35
cc_30 VNB N_VGND_c_387_n 0.0163916f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.725
cc_31 VNB N_VGND_c_388_n 0.0299087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_389_n 0.0164443f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.635
cc_33 VNB N_VGND_c_390_n 0.00629887f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.35
cc_34 VNB N_VGND_c_391_n 0.0107437f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.35
cc_35 VNB N_VGND_c_392_n 0.032693f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.71
cc_36 VNB N_VGND_c_393_n 0.0426063f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_37 VNB N_VGND_c_394_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.792 $Y2=1.685
cc_38 VNB N_VGND_c_395_n 0.230217f $X=-0.19 $Y=-0.245 $X2=1.792 $Y2=1.85
cc_39 VPB N_B_M1001_g 0.0514715f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_40 VPB N_B_M1006_g 0.0496702f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.725
cc_41 VPB N_B_c_74_n 0.00996319f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.565
cc_42 VPB N_B_c_76_n 0.0295401f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.35
cc_43 VPB B 0.00295203f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_44 VPB N_B_c_78_n 0.0208158f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.685
cc_45 VPB N_B_c_79_n 0.00371058f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.71
cc_46 VPB N_A_M1003_g 0.0185103f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_47 VPB N_A_M1000_g 0.0194047f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.725
cc_48 VPB N_A_c_156_n 0.0223344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_c_153_n 0.0319232f $X=-0.19 $Y=1.655 $X2=0.465 $Y2=1.35
cc_50 VPB N_A_27_481#_M1007_g 0.0279789f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=0.635
cc_51 VPB N_A_27_481#_c_214_n 0.0366122f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.35
cc_52 VPB N_A_27_481#_c_215_n 0.0350859f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.71
cc_53 VPB N_A_27_481#_c_216_n 0.0133386f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.71
cc_54 VPB N_A_27_481#_c_211_n 0.00751187f $X=-0.19 $Y=1.655 $X2=0.465 $Y2=1.69
cc_55 VPB N_VPWR_c_285_n 0.00565635f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.85
cc_56 VPB N_VPWR_c_286_n 0.00676633f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=1.52
cc_57 VPB N_VPWR_c_287_n 0.0275168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_288_n 0.00481431f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.565
cc_59 VPB N_VPWR_c_289_n 0.016633f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.35
cc_60 VPB N_VPWR_c_290_n 0.00430292f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.35
cc_61 VPB N_VPWR_c_291_n 0.0381457f $X=-0.19 $Y=1.655 $X2=0.465 $Y2=1.35
cc_62 VPB N_VPWR_c_284_n 0.0718012f $X=-0.19 $Y=1.655 $X2=0.465 $Y2=1.185
cc_63 VPB N_A_274_481#_c_323_n 0.00231305f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.85
cc_64 VPB N_A_274_481#_c_324_n 0.00715105f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.725
cc_65 VPB N_A_274_481#_c_325_n 0.00278331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_274_481#_c_326_n 0.0327489f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=1.52
cc_67 VPB N_A_274_481#_c_327_n 0.0466849f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.565
cc_68 VPB N_A_274_481#_c_328_n 0.0124855f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.35
cc_69 VPB N_X_c_357_n 0.00423602f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.635
cc_70 VPB N_X_c_358_n 0.00249605f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.85
cc_71 VPB N_X_c_355_n 0.00143791f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=1.52
cc_72 N_B_M1009_g N_A_M1002_g 0.0269706f $X=0.65 $Y=0.635 $X2=0 $Y2=0
cc_73 N_B_M1005_g N_A_M1004_g 0.0532399f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_74 N_B_M1001_g N_A_c_156_n 0.0552943f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_75 N_B_c_79_n N_A_c_156_n 0.00129594f $X=1.52 $Y=1.71 $X2=0 $Y2=0
cc_76 N_B_c_75_n N_A_c_151_n 2.06604e-19 $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_77 N_B_c_76_n N_A_c_151_n 0.0269706f $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_78 B N_A_c_151_n 0.00453346f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B_c_79_n N_A_c_151_n 0.00401433f $X=1.52 $Y=1.71 $X2=0 $Y2=0
cc_80 N_B_c_75_n A 0.0143205f $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_81 N_B_c_76_n A 0.0123935f $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_82 B A 0.0153065f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_83 N_B_c_79_n A 0.0537595f $X=1.52 $Y=1.71 $X2=0 $Y2=0
cc_84 N_B_M1001_g N_A_c_153_n 0.00752897f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_85 N_B_M1006_g N_A_c_153_n 0.0337099f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_86 N_B_M1005_g N_A_c_153_n 0.005063f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_87 N_B_c_75_n N_A_c_153_n 7.11439e-19 $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_88 B N_A_c_153_n 0.00605564f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B_c_78_n N_A_c_153_n 0.0180721f $X=1.775 $Y=1.685 $X2=0 $Y2=0
cc_90 N_B_c_79_n N_A_c_153_n 0.025605f $X=1.52 $Y=1.71 $X2=0 $Y2=0
cc_91 N_B_M1005_g N_A_27_481#_c_202_n 0.0172329f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_92 N_B_M1001_g N_A_27_481#_c_214_n 0.0194115f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_93 N_B_M1001_g N_A_27_481#_c_215_n 0.0112969f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_94 N_B_M1006_g N_A_27_481#_c_215_n 0.012315f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_95 N_B_c_74_n N_A_27_481#_c_215_n 0.00224846f $X=0.33 $Y=1.565 $X2=0 $Y2=0
cc_96 N_B_c_76_n N_A_27_481#_c_215_n 0.00460324f $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_97 B N_A_27_481#_c_215_n 0.0339094f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_98 N_B_c_78_n N_A_27_481#_c_215_n 0.00271895f $X=1.775 $Y=1.685 $X2=0 $Y2=0
cc_99 N_B_c_79_n N_A_27_481#_c_215_n 0.0792423f $X=1.52 $Y=1.71 $X2=0 $Y2=0
cc_100 N_B_M1001_g N_A_27_481#_c_216_n 0.00419608f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_101 N_B_c_74_n N_A_27_481#_c_216_n 0.0194805f $X=0.33 $Y=1.565 $X2=0 $Y2=0
cc_102 N_B_c_76_n N_A_27_481#_c_216_n 0.00152664f $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_103 N_B_M1009_g N_A_27_481#_c_206_n 0.00100576f $X=0.65 $Y=0.635 $X2=0 $Y2=0
cc_104 N_B_M1005_g N_A_27_481#_c_207_n 0.01618f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_105 B N_A_27_481#_c_207_n 0.0336809f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B_c_78_n N_A_27_481#_c_207_n 7.64722e-19 $X=1.775 $Y=1.685 $X2=0 $Y2=0
cc_107 N_B_c_79_n N_A_27_481#_c_207_n 0.00569422f $X=1.52 $Y=1.71 $X2=0 $Y2=0
cc_108 N_B_M1009_g N_A_27_481#_c_208_n 0.00572358f $X=0.65 $Y=0.635 $X2=0 $Y2=0
cc_109 N_B_M1005_g N_A_27_481#_c_209_n 0.00549818f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_110 B N_A_27_481#_c_209_n 0.0362021f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 B N_A_27_481#_c_210_n 4.9454e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B_c_78_n N_A_27_481#_c_210_n 0.0172329f $X=1.775 $Y=1.685 $X2=0 $Y2=0
cc_113 N_B_M1006_g N_A_27_481#_c_211_n 0.00454699f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_114 N_B_c_78_n N_A_27_481#_c_212_n 0.00549818f $X=1.775 $Y=1.685 $X2=0 $Y2=0
cc_115 N_B_M1001_g N_VPWR_c_285_n 0.00275065f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_116 N_B_M1006_g N_VPWR_c_286_n 0.00338591f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_117 N_B_M1001_g N_VPWR_c_287_n 0.00502664f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_118 N_B_M1006_g N_VPWR_c_289_n 0.0053602f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_119 N_B_M1001_g N_VPWR_c_284_n 0.0101321f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_120 N_B_M1006_g N_VPWR_c_284_n 0.00654225f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_121 N_B_M1006_g N_A_274_481#_c_324_n 0.0117414f $X=1.725 $Y=2.725 $X2=0 $Y2=0
cc_122 N_B_M1006_g N_A_274_481#_c_328_n 0.00322052f $X=1.725 $Y=2.725 $X2=0
+ $Y2=0
cc_123 N_B_M1005_g N_X_c_355_n 0.00288432f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_124 N_B_M1005_g N_X_c_356_n 0.00486523f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_125 N_B_M1009_g N_VGND_c_388_n 0.00395813f $X=0.65 $Y=0.635 $X2=0 $Y2=0
cc_126 N_B_c_75_n N_VGND_c_388_n 0.00855543f $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_127 N_B_c_76_n N_VGND_c_388_n 0.00454173f $X=0.37 $Y=1.35 $X2=0 $Y2=0
cc_128 N_B_M1009_g N_VGND_c_389_n 0.00537957f $X=0.65 $Y=0.635 $X2=0 $Y2=0
cc_129 N_B_M1009_g N_VGND_c_390_n 3.85551e-19 $X=0.65 $Y=0.635 $X2=0 $Y2=0
cc_130 N_B_M1005_g N_VGND_c_390_n 0.00140279f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_131 N_B_M1005_g N_VGND_c_393_n 0.00532993f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_132 N_B_M1009_g N_VGND_c_395_n 0.00528353f $X=0.65 $Y=0.635 $X2=0 $Y2=0
cc_133 N_B_M1005_g N_VGND_c_395_n 0.00528353f $X=1.9 $Y=0.635 $X2=0 $Y2=0
cc_134 N_A_c_156_n N_A_27_481#_c_214_n 0.00289801f $X=1.295 $Y=2.17 $X2=0 $Y2=0
cc_135 N_A_c_156_n N_A_27_481#_c_215_n 0.0271214f $X=1.295 $Y=2.17 $X2=0 $Y2=0
cc_136 N_A_c_153_n N_A_27_481#_c_215_n 0.00928444f $X=1.17 $Y=1.295 $X2=0 $Y2=0
cc_137 N_A_M1002_g N_A_27_481#_c_206_n 9.43578e-19 $X=1.08 $Y=0.635 $X2=0 $Y2=0
cc_138 N_A_M1002_g N_A_27_481#_c_207_n 0.0137683f $X=1.08 $Y=0.635 $X2=0 $Y2=0
cc_139 N_A_M1004_g N_A_27_481#_c_207_n 0.014244f $X=1.51 $Y=0.635 $X2=0 $Y2=0
cc_140 N_A_c_151_n N_A_27_481#_c_207_n 0.00289453f $X=1.51 $Y=1.205 $X2=0 $Y2=0
cc_141 A N_A_27_481#_c_207_n 0.0276411f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_142 A N_A_27_481#_c_208_n 0.0194543f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A_M1003_g N_VPWR_c_285_n 0.015859f $X=0.865 $Y=2.725 $X2=0 $Y2=0
cc_144 N_A_M1000_g N_VPWR_c_285_n 0.00172809f $X=1.295 $Y=2.725 $X2=0 $Y2=0
cc_145 N_A_c_156_n N_VPWR_c_285_n 0.00285785f $X=1.295 $Y=2.17 $X2=0 $Y2=0
cc_146 N_A_M1003_g N_VPWR_c_287_n 0.00445056f $X=0.865 $Y=2.725 $X2=0 $Y2=0
cc_147 N_A_M1000_g N_VPWR_c_289_n 0.0053602f $X=1.295 $Y=2.725 $X2=0 $Y2=0
cc_148 N_A_M1003_g N_VPWR_c_284_n 0.00804604f $X=0.865 $Y=2.725 $X2=0 $Y2=0
cc_149 N_A_M1000_g N_VPWR_c_284_n 0.0102021f $X=1.295 $Y=2.725 $X2=0 $Y2=0
cc_150 N_A_M1000_g N_A_274_481#_c_325_n 8.42648e-19 $X=1.295 $Y=2.725 $X2=0
+ $Y2=0
cc_151 N_A_M1004_g N_X_c_356_n 7.8665e-19 $X=1.51 $Y=0.635 $X2=0 $Y2=0
cc_152 N_A_M1002_g N_VGND_c_389_n 0.00447026f $X=1.08 $Y=0.635 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_VGND_c_390_n 0.00728733f $X=1.08 $Y=0.635 $X2=0 $Y2=0
cc_154 N_A_M1004_g N_VGND_c_390_n 0.00931849f $X=1.51 $Y=0.635 $X2=0 $Y2=0
cc_155 N_A_M1004_g N_VGND_c_393_n 0.00447026f $X=1.51 $Y=0.635 $X2=0 $Y2=0
cc_156 N_A_M1002_g N_VGND_c_395_n 0.00443817f $X=1.08 $Y=0.635 $X2=0 $Y2=0
cc_157 N_A_M1004_g N_VGND_c_395_n 0.00443817f $X=1.51 $Y=0.635 $X2=0 $Y2=0
cc_158 N_A_27_481#_c_214_n N_VPWR_c_285_n 0.0213595f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_159 N_A_27_481#_c_215_n N_VPWR_c_285_n 0.021643f $X=2.205 $Y=2.11 $X2=0 $Y2=0
cc_160 N_A_27_481#_c_214_n N_VPWR_c_287_n 0.0220321f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_161 N_A_27_481#_c_214_n N_VPWR_c_284_n 0.0125808f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_162 N_A_27_481#_c_215_n N_A_274_481#_c_324_n 0.0413416f $X=2.205 $Y=2.11
+ $X2=0 $Y2=0
cc_163 N_A_27_481#_c_215_n N_A_274_481#_c_325_n 0.0219276f $X=2.205 $Y=2.11
+ $X2=0 $Y2=0
cc_164 N_A_27_481#_M1007_g N_A_274_481#_c_326_n 0.00678379f $X=2.875 $Y=2.155
+ $X2=0 $Y2=0
cc_165 N_A_27_481#_M1007_g N_A_274_481#_c_327_n 0.00410645f $X=2.875 $Y=2.155
+ $X2=0 $Y2=0
cc_166 N_A_27_481#_M1007_g N_A_274_481#_c_328_n 0.00211575f $X=2.875 $Y=2.155
+ $X2=0 $Y2=0
cc_167 N_A_27_481#_c_215_n N_A_274_481#_c_328_n 0.015316f $X=2.205 $Y=2.11 $X2=0
+ $Y2=0
cc_168 N_A_27_481#_M1007_g N_X_c_357_n 0.00171503f $X=2.875 $Y=2.155 $X2=0 $Y2=0
cc_169 N_A_27_481#_c_211_n N_X_c_357_n 0.0160326f $X=2.29 $Y=2.025 $X2=0 $Y2=0
cc_170 N_A_27_481#_M1007_g N_X_c_358_n 0.00590235f $X=2.875 $Y=2.155 $X2=0 $Y2=0
cc_171 N_A_27_481#_c_215_n N_X_c_358_n 0.0145764f $X=2.205 $Y=2.11 $X2=0 $Y2=0
cc_172 N_A_27_481#_c_203_n N_X_c_354_n 0.00341197f $X=2.875 $Y=0.955 $X2=0 $Y2=0
cc_173 N_A_27_481#_c_201_n N_X_c_355_n 0.00919036f $X=2.8 $Y=1.03 $X2=0 $Y2=0
cc_174 N_A_27_481#_c_203_n N_X_c_355_n 0.0100263f $X=2.875 $Y=0.955 $X2=0 $Y2=0
cc_175 N_A_27_481#_M1007_g N_X_c_355_n 0.0348859f $X=2.875 $Y=2.155 $X2=0 $Y2=0
cc_176 N_A_27_481#_c_205_n N_X_c_355_n 0.00593165f $X=2.875 $Y=1.03 $X2=0 $Y2=0
cc_177 N_A_27_481#_c_207_n N_X_c_355_n 0.0136536f $X=2.205 $Y=0.955 $X2=0 $Y2=0
cc_178 N_A_27_481#_c_209_n N_X_c_355_n 0.042946f $X=2.38 $Y=1.12 $X2=0 $Y2=0
cc_179 N_A_27_481#_c_210_n N_X_c_355_n 0.0035089f $X=2.38 $Y=1.12 $X2=0 $Y2=0
cc_180 N_A_27_481#_c_211_n N_X_c_355_n 0.0103172f $X=2.29 $Y=2.025 $X2=0 $Y2=0
cc_181 N_A_27_481#_c_202_n N_X_c_356_n 0.0081728f $X=2.545 $Y=1.03 $X2=0 $Y2=0
cc_182 N_A_27_481#_c_207_n N_X_c_356_n 0.0390086f $X=2.205 $Y=0.955 $X2=0 $Y2=0
cc_183 N_A_27_481#_c_206_n N_VGND_c_388_n 0.00232547f $X=0.865 $Y=0.635 $X2=0
+ $Y2=0
cc_184 N_A_27_481#_c_206_n N_VGND_c_389_n 0.00857925f $X=0.865 $Y=0.635 $X2=0
+ $Y2=0
cc_185 N_A_27_481#_c_206_n N_VGND_c_390_n 0.0125867f $X=0.865 $Y=0.635 $X2=0
+ $Y2=0
cc_186 N_A_27_481#_c_207_n N_VGND_c_390_n 0.0216087f $X=2.205 $Y=0.955 $X2=0
+ $Y2=0
cc_187 N_A_27_481#_c_203_n N_VGND_c_392_n 0.005455f $X=2.875 $Y=0.955 $X2=0
+ $Y2=0
cc_188 N_A_27_481#_c_203_n N_VGND_c_393_n 0.00523054f $X=2.875 $Y=0.955 $X2=0
+ $Y2=0
cc_189 N_A_27_481#_c_203_n N_VGND_c_395_n 0.00528353f $X=2.875 $Y=0.955 $X2=0
+ $Y2=0
cc_190 N_A_27_481#_c_206_n N_VGND_c_395_n 0.00817244f $X=0.865 $Y=0.635 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_285_n N_A_274_481#_c_323_n 0.00153963f $X=1.08 $Y=2.55 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_286_n N_A_274_481#_c_323_n 0.00150838f $X=1.94 $Y=2.87 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_289_n N_A_274_481#_c_323_n 0.0173997f $X=1.81 $Y=3.33 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_284_n N_A_274_481#_c_323_n 0.0099853f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_VPWR_M1006_d N_A_274_481#_c_324_n 0.00305508f $X=1.8 $Y=2.405 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_286_n N_A_274_481#_c_324_n 0.0140774f $X=1.94 $Y=2.87 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_284_n N_A_274_481#_c_324_n 0.0119298f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_285_n N_A_274_481#_c_325_n 0.00166618f $X=1.08 $Y=2.55 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_291_n N_A_274_481#_c_326_n 0.0230291f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_284_n N_A_274_481#_c_326_n 0.0284686f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_286_n N_A_274_481#_c_328_n 0.00981802f $X=1.94 $Y=2.87 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_291_n N_A_274_481#_c_328_n 0.0045837f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_284_n N_A_274_481#_c_328_n 0.00555566f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_204 N_A_274_481#_c_327_n N_X_c_357_n 0.02624f $X=3.09 $Y=1.98 $X2=0 $Y2=0
cc_205 N_A_274_481#_c_326_n N_X_c_358_n 0.0219496f $X=2.985 $Y=2.75 $X2=0 $Y2=0
cc_206 N_A_274_481#_c_328_n N_X_c_358_n 0.0099835f $X=2.29 $Y=2.45 $X2=0 $Y2=0
cc_207 N_X_c_356_n N_VGND_c_390_n 0.00934303f $X=2.645 $Y=0.555 $X2=0 $Y2=0
cc_208 N_X_c_354_n N_VGND_c_392_n 0.0127834f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_209 N_X_c_354_n N_VGND_c_393_n 0.00606568f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_210 N_X_c_356_n N_VGND_c_393_n 0.0227309f $X=2.645 $Y=0.555 $X2=0 $Y2=0
cc_211 N_X_c_354_n N_VGND_c_395_n 0.0060325f $X=2.73 $Y=0.7 $X2=0 $Y2=0
cc_212 N_X_c_356_n N_VGND_c_395_n 0.0232607f $X=2.645 $Y=0.555 $X2=0 $Y2=0
