* File: sky130_fd_sc_lp__mux2_4.spice
* Created: Fri Aug 28 10:44:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2_4.pex.spice"
.subckt sky130_fd_sc_lp__mux2_4  VNB VPB S A0 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_S_M1007_g N_A_41_367#_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1722 AS=0.2226 PD=1.25 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1008 A_287_47# N_A_41_367#_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1722 PD=1.05 PS=1.25 NRD=7.14 NRS=9.276 M=1 R=5.6 SA=75000.7
+ SB=75003.8 A=0.126 P=1.98 MULT=1
MM1010 N_A_359_47#_M1010_d N_A0_M1010_g A_287_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2499 AS=0.0882 PD=1.435 PS=1.05 NRD=44.988 NRS=7.14 M=1 R=5.6 SA=75001.1
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1011 A_508_47# N_A1_M1011_g N_A_359_47#_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2499 PD=1.05 PS=1.435 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_S_M1004_g A_508_47# VNB NSHORT L=0.15 W=0.84 AD=0.2898
+ AS=0.0882 PD=1.53 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75002.2 SB=75002.3
+ A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1004_d N_A_359_47#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2898 AS=0.1176 PD=1.53 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A_359_47#_M1001_g N_X_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1001_d N_A_359_47#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_A_359_47#_M1015_g N_X_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_S_M1013_g N_A_41_367#_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_A_210_367#_M1017_d N_A_41_367#_M1017_g N_VPWR_M1013_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_359_47#_M1005_d N_A0_M1005_g N_A_317_367#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1002 N_A_210_367#_M1002_d N_A1_M1002_g N_A_359_47#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_S_M1009_g N_A_317_367#_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_X_M1003_d N_A_359_47#_M1003_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_X_M1003_d N_A_359_47#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1012 N_X_M1012_d N_A_359_47#_M1012_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_X_M1012_d N_A_359_47#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__mux2_4.pxi.spice"
*
.ends
*
*
