# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__decapkapwr_8
  CLASS CORE SPACER ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__decapkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.495000 2.105000 0.905000 2.675000 ;
        RECT 0.495000 2.675000 3.285000 2.945000 ;
        RECT 0.495000 2.945000 0.905000 3.075000 ;
        RECT 1.955000 1.340000 3.285000 1.675000 ;
        RECT 2.865000 1.675000 3.285000 2.675000 ;
        RECT 2.865000 2.945000 3.285000 3.075000 ;
      LAYER mcon ;
        RECT 0.575000 2.725000 0.745000 2.895000 ;
        RECT 0.940000 2.725000 1.110000 2.895000 ;
        RECT 1.345000 2.725000 1.515000 2.895000 ;
        RECT 1.765000 2.725000 1.935000 2.895000 ;
        RECT 2.170000 2.725000 2.340000 2.895000 ;
        RECT 2.565000 2.725000 2.735000 2.895000 ;
        RECT 3.025000 2.725000 3.195000 2.895000 ;
      LAYER met1 ;
        RECT 0.070000 2.675000 3.770000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
        RECT 0.650000  0.085000 0.980000 1.605000 ;
        RECT 0.650000  1.605000 1.560000 1.935000 ;
        RECT 2.930000  0.085000 3.260000 1.125000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.840000 3.415000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
END sky130_fd_sc_lp__decapkapwr_8
