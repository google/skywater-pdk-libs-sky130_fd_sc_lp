* File: sky130_fd_sc_lp__o21ai_m.spice
* Created: Fri Aug 28 11:05:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o21ai_m  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_27_51#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_27_51#_M1000_d N_A2_M1000_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_27_51#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_110_434# N_A1_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A2_M1003_g A_110_434# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=51.5943 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
c_24 VNB 0 1.57953e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o21ai_m.pxi.spice"
*
.ends
*
*
