* File: sky130_fd_sc_lp__a31oi_2.pxi.spice
* Created: Fri Aug 28 10:00:05 2020
* 
x_PM_SKY130_FD_SC_LP__A31OI_2%A3 N_A3_c_81_n N_A3_M1009_g N_A3_M1005_g
+ N_A3_c_83_n N_A3_c_84_n N_A3_M1012_g N_A3_M1014_g N_A3_c_86_n A3 N_A3_c_88_n
+ PM_SKY130_FD_SC_LP__A31OI_2%A3
x_PM_SKY130_FD_SC_LP__A31OI_2%A2 N_A2_c_128_n N_A2_M1003_g N_A2_M1000_g
+ N_A2_c_130_n N_A2_M1011_g N_A2_M1001_g A2 A2 N_A2_c_132_n N_A2_c_133_n
+ PM_SKY130_FD_SC_LP__A31OI_2%A2
x_PM_SKY130_FD_SC_LP__A31OI_2%A1 N_A1_M1002_g N_A1_c_185_n N_A1_c_186_n
+ N_A1_M1007_g N_A1_c_188_n N_A1_M1015_g N_A1_M1008_g N_A1_c_190_n A1
+ N_A1_c_191_n N_A1_c_192_n PM_SKY130_FD_SC_LP__A31OI_2%A1
x_PM_SKY130_FD_SC_LP__A31OI_2%B1 N_B1_M1006_g N_B1_M1004_g N_B1_M1013_g
+ N_B1_M1010_g B1 B1 B1 N_B1_c_253_n PM_SKY130_FD_SC_LP__A31OI_2%B1
x_PM_SKY130_FD_SC_LP__A31OI_2%A_27_367# N_A_27_367#_M1005_d N_A_27_367#_M1014_d
+ N_A_27_367#_M1001_s N_A_27_367#_M1008_d N_A_27_367#_M1010_d
+ N_A_27_367#_c_294_n N_A_27_367#_c_295_n N_A_27_367#_c_296_n
+ N_A_27_367#_c_326_p N_A_27_367#_c_297_n N_A_27_367#_c_316_n
+ N_A_27_367#_c_348_p N_A_27_367#_c_318_n N_A_27_367#_c_329_p
+ N_A_27_367#_c_298_n N_A_27_367#_c_299_n N_A_27_367#_c_300_n
+ N_A_27_367#_c_342_p PM_SKY130_FD_SC_LP__A31OI_2%A_27_367#
x_PM_SKY130_FD_SC_LP__A31OI_2%VPWR N_VPWR_M1005_s N_VPWR_M1000_d N_VPWR_M1002_s
+ N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n VPWR
+ N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_355_n N_VPWR_c_363_n N_VPWR_c_364_n
+ N_VPWR_c_365_n PM_SKY130_FD_SC_LP__A31OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A31OI_2%Y N_Y_M1007_s N_Y_M1015_s N_Y_M1013_s N_Y_M1004_s
+ N_Y_c_419_n N_Y_c_420_n N_Y_c_438_n N_Y_c_421_n N_Y_c_422_n N_Y_c_423_n
+ N_Y_c_424_n N_Y_c_425_n N_Y_c_444_n Y Y PM_SKY130_FD_SC_LP__A31OI_2%Y
x_PM_SKY130_FD_SC_LP__A31OI_2%A_27_69# N_A_27_69#_M1009_s N_A_27_69#_M1012_s
+ N_A_27_69#_M1011_s N_A_27_69#_c_495_n N_A_27_69#_c_496_n N_A_27_69#_c_502_n
+ N_A_27_69#_c_497_n N_A_27_69#_c_509_n N_A_27_69#_c_513_n N_A_27_69#_c_498_n
+ PM_SKY130_FD_SC_LP__A31OI_2%A_27_69#
x_PM_SKY130_FD_SC_LP__A31OI_2%VGND N_VGND_M1009_d N_VGND_M1006_d N_VGND_c_537_n
+ N_VGND_c_538_n N_VGND_c_539_n N_VGND_c_540_n VGND N_VGND_c_541_n
+ N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n PM_SKY130_FD_SC_LP__A31OI_2%VGND
x_PM_SKY130_FD_SC_LP__A31OI_2%A_282_69# N_A_282_69#_M1003_d N_A_282_69#_M1007_d
+ N_A_282_69#_c_589_n N_A_282_69#_c_595_n N_A_282_69#_c_590_n
+ PM_SKY130_FD_SC_LP__A31OI_2%A_282_69#
cc_1 VNB N_A3_c_81_n 0.0213789f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_2 VNB N_A3_M1005_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A3_c_83_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.37
cc_4 VNB N_A3_c_84_n 0.0159218f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.295
cc_5 VNB N_A3_M1014_g 0.0100053f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_6 VNB N_A3_c_86_n 0.00438315f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.37
cc_7 VNB A3 0.0157429f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A3_c_88_n 0.0435904f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.46
cc_9 VNB N_A2_c_128_n 0.0164944f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_10 VNB N_A2_M1000_g 0.00161519f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_11 VNB N_A2_c_130_n 0.0196299f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.37
cc_12 VNB N_A2_M1001_g 0.001613f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.445
cc_13 VNB N_A2_c_132_n 0.0130901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_133_n 0.0443925f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.46
cc_15 VNB N_A1_M1002_g 0.00925787f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_16 VNB N_A1_c_185_n 0.021447f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_17 VNB N_A1_c_186_n 0.013308f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_18 VNB N_A1_M1007_g 0.0232887f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.37
cc_19 VNB N_A1_c_188_n 0.0120334f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.765
cc_20 VNB N_A1_M1015_g 0.0196655f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_21 VNB N_A1_c_190_n 0.00665797f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_22 VNB N_A1_c_191_n 0.0223119f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_23 VNB N_A1_c_192_n 0.00122154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_M1006_g 0.0186619f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_25 VNB N_B1_M1013_g 0.0250995f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.765
cc_26 VNB B1 0.0267334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_c_253_n 0.0365303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_355_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_419_n 0.00460399f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_30 VNB N_Y_c_420_n 0.00569895f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.37
cc_31 VNB N_Y_c_421_n 0.00189149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_422_n 0.0128634f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.46
cc_33 VNB N_Y_c_423_n 0.0309544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_424_n 0.00178269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_425_n 0.00679811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.00223048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_69#_c_495_n 0.00751114f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.295
cc_38 VNB N_A_27_69#_c_496_n 0.0222114f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.765
cc_39 VNB N_A_27_69#_c_497_n 0.00209149f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_40 VNB N_A_27_69#_c_498_n 0.00982722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_537_n 0.00332106f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.37
cc_42 VNB N_VGND_c_538_n 0.00332106f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.445
cc_43 VNB N_VGND_c_539_n 0.0697434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_540_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.37
cc_45 VNB N_VGND_c_541_n 0.0165321f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_46 VNB N_VGND_c_542_n 0.0240479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_543_n 0.285644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_544_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_282_69#_c_589_n 0.018507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_282_69#_c_590_n 0.00278584f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.445
cc_51 VPB N_A3_M1005_g 0.0248454f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_52 VPB N_A3_M1014_g 0.0187449f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_53 VPB N_A2_M1000_g 0.0198852f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_54 VPB N_A2_M1001_g 0.0198864f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.445
cc_55 VPB N_A1_M1002_g 0.0238132f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_56 VPB N_A1_M1008_g 0.0219448f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A1_c_191_n 0.00663614f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.46
cc_58 VPB N_A1_c_192_n 0.00338102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B1_M1004_g 0.0183424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_B1_M1010_g 0.0244533f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_61 VPB B1 0.0226422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_B1_c_253_n 0.00489715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_27_367#_c_294_n 0.0450352f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_64 VPB N_A_27_367#_c_295_n 0.00352183f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_65 VPB N_A_27_367#_c_296_n 0.00915646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_27_367#_c_297_n 0.0087208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_27_367#_c_298_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_27_367#_c_299_n 0.0374018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_27_367#_c_300_n 0.00220677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_356_n 4.06898e-19 $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.765
cc_71 VPB N_VPWR_c_357_n 0.00431911f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_72 VPB N_VPWR_c_358_n 0.0149824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_359_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.46
cc_74 VPB N_VPWR_c_360_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_361_n 0.0419995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_355_n 0.0548462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_363_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_364_n 0.0147652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_365_n 0.0167608f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB Y 0.00324587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 N_A3_c_84_n N_A2_c_128_n 0.0174534f $X=0.905 $Y=1.295 $X2=-0.19 $Y2=-0.245
cc_82 N_A3_M1014_g N_A2_M1000_g 0.0174534f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A3_c_81_n N_A2_c_132_n 6.46746e-19 $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_84 N_A3_c_83_n N_A2_c_132_n 0.00826423f $X=0.83 $Y=1.37 $X2=0 $Y2=0
cc_85 N_A3_c_84_n N_A2_c_132_n 0.00497493f $X=0.905 $Y=1.295 $X2=0 $Y2=0
cc_86 N_A3_M1014_g N_A2_c_132_n 0.00549183f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A3_c_86_n N_A2_c_132_n 0.00391242f $X=0.905 $Y=1.37 $X2=0 $Y2=0
cc_88 A3 N_A2_c_132_n 0.0275616f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A3_c_88_n N_A2_c_132_n 8.74451e-19 $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_90 N_A3_c_86_n N_A2_c_133_n 0.0174534f $X=0.905 $Y=1.37 $X2=0 $Y2=0
cc_91 N_A3_M1005_g N_A_27_367#_c_295_n 0.0161348f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A3_c_83_n N_A_27_367#_c_295_n 5.52567e-19 $X=0.83 $Y=1.37 $X2=0 $Y2=0
cc_93 N_A3_M1014_g N_A_27_367#_c_295_n 0.013661f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_94 A3 N_A_27_367#_c_295_n 0.00724563f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_95 N_A3_c_88_n N_A_27_367#_c_295_n 0.00110593f $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_96 A3 N_A_27_367#_c_296_n 0.0221781f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A3_c_88_n N_A_27_367#_c_296_n 0.00590098f $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_98 N_A3_M1005_g N_VPWR_c_356_n 0.0169864f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A3_M1014_g N_VPWR_c_356_n 0.0150873f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A3_M1014_g N_VPWR_c_358_n 0.00486043f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A3_M1005_g N_VPWR_c_360_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A3_M1005_g N_VPWR_c_355_n 0.00917987f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A3_M1014_g N_VPWR_c_355_n 0.0082726f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_104 A3 N_A_27_69#_c_495_n 0.0218403f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A3_c_88_n N_A_27_69#_c_495_n 0.00139244f $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_106 N_A3_c_81_n N_A_27_69#_c_496_n 0.00146542f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_107 N_A3_c_81_n N_A_27_69#_c_502_n 0.0135475f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_108 N_A3_c_83_n N_A_27_69#_c_502_n 5.72217e-19 $X=0.83 $Y=1.37 $X2=0 $Y2=0
cc_109 N_A3_c_84_n N_A_27_69#_c_502_n 0.012081f $X=0.905 $Y=1.295 $X2=0 $Y2=0
cc_110 A3 N_A_27_69#_c_502_n 0.00615389f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A3_c_84_n N_A_27_69#_c_497_n 3.49657e-19 $X=0.905 $Y=1.295 $X2=0 $Y2=0
cc_112 N_A3_c_81_n N_VGND_c_537_n 0.0113295f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_113 N_A3_c_84_n N_VGND_c_537_n 0.00876445f $X=0.905 $Y=1.295 $X2=0 $Y2=0
cc_114 N_A3_c_84_n N_VGND_c_539_n 0.00400407f $X=0.905 $Y=1.295 $X2=0 $Y2=0
cc_115 N_A3_c_81_n N_VGND_c_541_n 0.00400407f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_116 N_A3_c_81_n N_VGND_c_543_n 0.00796025f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_117 N_A3_c_84_n N_VGND_c_543_n 0.00775088f $X=0.905 $Y=1.295 $X2=0 $Y2=0
cc_118 N_A2_M1001_g N_A1_M1002_g 0.017836f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A2_c_132_n N_A1_c_186_n 8.31481e-19 $X=1.47 $Y=1.46 $X2=0 $Y2=0
cc_120 N_A2_c_133_n N_A1_c_186_n 0.017836f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_121 N_A2_c_132_n N_A_27_367#_c_295_n 0.0305315f $X=1.47 $Y=1.46 $X2=0 $Y2=0
cc_122 N_A2_M1000_g N_A_27_367#_c_297_n 0.0134371f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A2_M1001_g N_A_27_367#_c_297_n 0.0161877f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A2_c_132_n N_A_27_367#_c_297_n 0.0276211f $X=1.47 $Y=1.46 $X2=0 $Y2=0
cc_125 N_A2_c_133_n N_A_27_367#_c_297_n 0.00503764f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_126 N_A2_M1000_g N_A_27_367#_c_300_n 0.00138835f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_A2_c_132_n N_A_27_367#_c_300_n 0.0208108f $X=1.47 $Y=1.46 $X2=0 $Y2=0
cc_128 N_A2_M1000_g N_VPWR_c_356_n 7.56711e-19 $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A2_M1000_g N_VPWR_c_357_n 0.00188227f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A2_M1001_g N_VPWR_c_357_n 0.00191629f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A2_M1000_g N_VPWR_c_358_n 0.00585385f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A2_M1000_g N_VPWR_c_355_n 0.0107688f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A2_M1001_g N_VPWR_c_355_n 0.0107415f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A2_M1001_g N_VPWR_c_364_n 0.00585385f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A2_M1001_g N_VPWR_c_365_n 6.04823e-19 $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_c_130_n N_Y_c_424_n 0.00173106f $X=1.765 $Y=1.295 $X2=0 $Y2=0
cc_137 N_A2_c_130_n Y 0.00107159f $X=1.765 $Y=1.295 $X2=0 $Y2=0
cc_138 N_A2_c_133_n Y 0.00375305f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_139 N_A2_c_132_n N_A_27_69#_c_502_n 0.0264982f $X=1.47 $Y=1.46 $X2=0 $Y2=0
cc_140 N_A2_c_128_n N_A_27_69#_c_497_n 3.80426e-19 $X=1.335 $Y=1.295 $X2=0 $Y2=0
cc_141 N_A2_c_128_n N_A_27_69#_c_509_n 0.0127808f $X=1.335 $Y=1.295 $X2=0 $Y2=0
cc_142 N_A2_c_130_n N_A_27_69#_c_509_n 0.011004f $X=1.765 $Y=1.295 $X2=0 $Y2=0
cc_143 N_A2_c_132_n N_A_27_69#_c_509_n 0.0263173f $X=1.47 $Y=1.46 $X2=0 $Y2=0
cc_144 N_A2_c_133_n N_A_27_69#_c_509_n 5.64665e-19 $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_145 N_A2_c_132_n N_A_27_69#_c_513_n 0.0171283f $X=1.47 $Y=1.46 $X2=0 $Y2=0
cc_146 N_A2_c_128_n N_A_27_69#_c_498_n 0.00135967f $X=1.335 $Y=1.295 $X2=0 $Y2=0
cc_147 N_A2_c_130_n N_A_27_69#_c_498_n 0.00926257f $X=1.765 $Y=1.295 $X2=0 $Y2=0
cc_148 N_A2_c_133_n N_A_27_69#_c_498_n 0.0028277f $X=1.845 $Y=1.46 $X2=0 $Y2=0
cc_149 N_A2_c_128_n N_VGND_c_537_n 6.22792e-19 $X=1.335 $Y=1.295 $X2=0 $Y2=0
cc_150 N_A2_c_128_n N_VGND_c_539_n 0.00482246f $X=1.335 $Y=1.295 $X2=0 $Y2=0
cc_151 N_A2_c_130_n N_VGND_c_539_n 0.0029147f $X=1.765 $Y=1.295 $X2=0 $Y2=0
cc_152 N_A2_c_128_n N_VGND_c_543_n 0.00955107f $X=1.335 $Y=1.295 $X2=0 $Y2=0
cc_153 N_A2_c_130_n N_VGND_c_543_n 0.00428625f $X=1.765 $Y=1.295 $X2=0 $Y2=0
cc_154 N_A2_c_130_n N_A_282_69#_c_589_n 0.0112238f $X=1.765 $Y=1.295 $X2=0 $Y2=0
cc_155 N_A2_c_128_n N_A_282_69#_c_590_n 0.00115849f $X=1.335 $Y=1.295 $X2=0
+ $Y2=0
cc_156 N_A1_M1015_g N_B1_M1006_g 0.018756f $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_157 N_A1_M1008_g N_B1_M1004_g 0.036457f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A1_c_192_n N_B1_M1004_g 2.20954e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A1_M1008_g B1 2.72793e-19 $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A1_c_191_n B1 0.00169089f $X=3.17 $Y=1.42 $X2=0 $Y2=0
cc_161 N_A1_c_192_n B1 0.027789f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A1_c_191_n N_B1_c_253_n 0.0188144f $X=3.17 $Y=1.42 $X2=0 $Y2=0
cc_163 N_A1_c_192_n N_B1_c_253_n 2.70573e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A1_M1002_g N_A_27_367#_c_297_n 0.00100697f $X=2.275 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A1_M1002_g N_A_27_367#_c_316_n 0.0158963f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A1_M1008_g N_A_27_367#_c_316_n 0.011818f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A1_M1008_g N_VPWR_c_361_n 0.00486043f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A1_M1002_g N_VPWR_c_355_n 0.00458845f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A1_M1008_g N_VPWR_c_355_n 0.00458845f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A1_M1002_g N_VPWR_c_364_n 0.00486043f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A1_M1002_g N_VPWR_c_365_n 0.013564f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A1_M1008_g N_VPWR_c_365_n 0.0146909f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A1_M1007_g N_Y_c_419_n 0.00711362f $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_174 N_A1_M1015_g N_Y_c_419_n 2.76958e-19 $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_175 N_A1_M1007_g N_Y_c_420_n 0.00248848f $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_176 N_A1_c_188_n N_Y_c_420_n 0.00509897f $X=3.005 $Y=1.42 $X2=0 $Y2=0
cc_177 N_A1_M1015_g N_Y_c_420_n 0.0134854f $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_178 N_A1_c_191_n N_Y_c_420_n 8.78513e-19 $X=3.17 $Y=1.42 $X2=0 $Y2=0
cc_179 N_A1_c_192_n N_Y_c_420_n 0.0275407f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A1_M1008_g N_Y_c_438_n 0.0131718f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A1_c_190_n N_Y_c_438_n 0.00484624f $X=2.72 $Y=1.42 $X2=0 $Y2=0
cc_182 N_A1_c_191_n N_Y_c_438_n 7.00572e-19 $X=3.17 $Y=1.42 $X2=0 $Y2=0
cc_183 N_A1_c_192_n N_Y_c_438_n 0.022079f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A1_M1015_g N_Y_c_421_n 8.28478e-19 $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_185 N_A1_M1007_g N_Y_c_424_n 0.00719778f $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_186 N_A1_M1008_g N_Y_c_444_n 7.61713e-19 $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A1_M1002_g Y 0.0154749f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A1_c_185_n Y 0.0180754f $X=2.645 $Y=1.42 $X2=0 $Y2=0
cc_189 N_A1_c_186_n Y 0.00308813f $X=2.35 $Y=1.42 $X2=0 $Y2=0
cc_190 N_A1_M1007_g Y 0.00433237f $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_191 N_A1_M1015_g Y 5.17418e-19 $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_192 N_A1_M1008_g Y 0.00666541f $X=3.225 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A1_c_190_n Y 0.0101725f $X=2.72 $Y=1.42 $X2=0 $Y2=0
cc_194 N_A1_c_191_n Y 7.4938e-19 $X=3.17 $Y=1.42 $X2=0 $Y2=0
cc_195 N_A1_c_192_n Y 0.0274037f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A1_M1002_g Y 0.00625946f $X=2.275 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A1_M1007_g N_A_27_69#_c_498_n 9.70779e-19 $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_198 N_A1_M1015_g N_VGND_c_538_n 6.53017e-19 $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_199 N_A1_M1007_g N_VGND_c_539_n 0.0029147f $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_200 N_A1_M1015_g N_VGND_c_539_n 0.00450424f $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_201 N_A1_M1007_g N_VGND_c_543_n 0.00432836f $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_202 N_A1_M1015_g N_VGND_c_543_n 0.00866668f $X=3.225 $Y=0.765 $X2=0 $Y2=0
cc_203 N_A1_M1007_g N_A_282_69#_c_589_n 0.0140502f $X=2.72 $Y=0.765 $X2=0 $Y2=0
cc_204 N_A1_M1015_g N_A_282_69#_c_589_n 0.00377143f $X=3.225 $Y=0.765 $X2=0
+ $Y2=0
cc_205 N_A1_M1015_g N_A_282_69#_c_595_n 0.00517317f $X=3.225 $Y=0.765 $X2=0
+ $Y2=0
cc_206 N_B1_M1004_g N_A_27_367#_c_318_n 0.0115031f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B1_M1010_g N_A_27_367#_c_318_n 0.0114565f $X=4.085 $Y=2.465 $X2=0 $Y2=0
cc_208 B1 N_A_27_367#_c_299_n 0.0219167f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_209 N_B1_M1004_g N_VPWR_c_361_n 0.00357877f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B1_M1010_g N_VPWR_c_361_n 0.00357877f $X=4.085 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B1_M1004_g N_VPWR_c_355_n 0.00537654f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_212 N_B1_M1010_g N_VPWR_c_355_n 0.00644538f $X=4.085 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B1_M1004_g N_VPWR_c_365_n 0.00116005f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_214 N_B1_M1004_g N_Y_c_438_n 0.0115282f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_215 B1 N_Y_c_438_n 0.011195f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_216 N_B1_M1006_g N_Y_c_421_n 8.28776e-19 $X=3.655 $Y=0.765 $X2=0 $Y2=0
cc_217 N_B1_M1006_g N_Y_c_422_n 0.013073f $X=3.655 $Y=0.765 $X2=0 $Y2=0
cc_218 N_B1_M1013_g N_Y_c_422_n 0.0136535f $X=4.085 $Y=0.765 $X2=0 $Y2=0
cc_219 B1 N_Y_c_422_n 0.0724456f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B1_c_253_n N_Y_c_422_n 0.00246472f $X=4.085 $Y=1.51 $X2=0 $Y2=0
cc_221 N_B1_M1013_g N_Y_c_423_n 0.00354556f $X=4.085 $Y=0.765 $X2=0 $Y2=0
cc_222 B1 N_Y_c_425_n 0.00265095f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_223 N_B1_M1004_g N_Y_c_444_n 0.0104433f $X=3.655 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B1_M1010_g N_Y_c_444_n 0.0109326f $X=4.085 $Y=2.465 $X2=0 $Y2=0
cc_225 B1 N_Y_c_444_n 0.0204377f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_226 N_B1_c_253_n N_Y_c_444_n 6.50093e-19 $X=4.085 $Y=1.51 $X2=0 $Y2=0
cc_227 N_B1_M1006_g N_VGND_c_538_n 0.0103777f $X=3.655 $Y=0.765 $X2=0 $Y2=0
cc_228 N_B1_M1013_g N_VGND_c_538_n 0.0127653f $X=4.085 $Y=0.765 $X2=0 $Y2=0
cc_229 N_B1_M1006_g N_VGND_c_539_n 0.00400407f $X=3.655 $Y=0.765 $X2=0 $Y2=0
cc_230 N_B1_M1013_g N_VGND_c_542_n 0.00400407f $X=4.085 $Y=0.765 $X2=0 $Y2=0
cc_231 N_B1_M1006_g N_VGND_c_543_n 0.00775088f $X=3.655 $Y=0.765 $X2=0 $Y2=0
cc_232 N_B1_M1013_g N_VGND_c_543_n 0.00799754f $X=4.085 $Y=0.765 $X2=0 $Y2=0
cc_233 N_B1_M1006_g N_A_282_69#_c_589_n 2.3575e-19 $X=3.655 $Y=0.765 $X2=0 $Y2=0
cc_234 N_A_27_367#_c_295_n N_VPWR_M1005_s 0.00176461f $X=1.025 $Y=1.8 $X2=-0.19
+ $Y2=1.655
cc_235 N_A_27_367#_c_297_n N_VPWR_M1000_d 0.00261503f $X=1.93 $Y=1.8 $X2=0 $Y2=0
cc_236 N_A_27_367#_c_316_n N_VPWR_M1002_s 0.018527f $X=3.345 $Y=2.385 $X2=0
+ $Y2=0
cc_237 N_A_27_367#_c_295_n N_VPWR_c_356_n 0.0170777f $X=1.025 $Y=1.8 $X2=0 $Y2=0
cc_238 N_A_27_367#_c_297_n N_VPWR_c_357_n 0.0200142f $X=1.93 $Y=1.8 $X2=0 $Y2=0
cc_239 N_A_27_367#_c_326_p N_VPWR_c_358_n 0.0140491f $X=1.12 $Y=1.98 $X2=0 $Y2=0
cc_240 N_A_27_367#_c_294_n N_VPWR_c_360_n 0.0178111f $X=0.26 $Y=1.98 $X2=0 $Y2=0
cc_241 N_A_27_367#_c_318_n N_VPWR_c_361_n 0.0361172f $X=4.205 $Y=2.99 $X2=0
+ $Y2=0
cc_242 N_A_27_367#_c_329_p N_VPWR_c_361_n 0.0125234f $X=3.535 $Y=2.99 $X2=0
+ $Y2=0
cc_243 N_A_27_367#_c_298_n N_VPWR_c_361_n 0.0179183f $X=4.335 $Y=2.905 $X2=0
+ $Y2=0
cc_244 N_A_27_367#_M1005_d N_VPWR_c_355_n 0.00371702f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_245 N_A_27_367#_M1014_d N_VPWR_c_355_n 0.00380103f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_246 N_A_27_367#_M1001_s N_VPWR_c_355_n 0.00288026f $X=1.92 $Y=1.835 $X2=0
+ $Y2=0
cc_247 N_A_27_367#_M1008_d N_VPWR_c_355_n 0.00254061f $X=3.3 $Y=1.835 $X2=0
+ $Y2=0
cc_248 N_A_27_367#_M1010_d N_VPWR_c_355_n 0.00215161f $X=4.16 $Y=1.835 $X2=0
+ $Y2=0
cc_249 N_A_27_367#_c_294_n N_VPWR_c_355_n 0.0100304f $X=0.26 $Y=1.98 $X2=0 $Y2=0
cc_250 N_A_27_367#_c_326_p N_VPWR_c_355_n 0.0090585f $X=1.12 $Y=1.98 $X2=0 $Y2=0
cc_251 N_A_27_367#_c_316_n N_VPWR_c_355_n 0.0119101f $X=3.345 $Y=2.385 $X2=0
+ $Y2=0
cc_252 N_A_27_367#_c_318_n N_VPWR_c_355_n 0.023676f $X=4.205 $Y=2.99 $X2=0 $Y2=0
cc_253 N_A_27_367#_c_329_p N_VPWR_c_355_n 0.0073762f $X=3.535 $Y=2.99 $X2=0
+ $Y2=0
cc_254 N_A_27_367#_c_298_n N_VPWR_c_355_n 0.0101029f $X=4.335 $Y=2.905 $X2=0
+ $Y2=0
cc_255 N_A_27_367#_c_342_p N_VPWR_c_355_n 0.00905721f $X=2.06 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_A_27_367#_c_342_p N_VPWR_c_364_n 0.0136943f $X=2.06 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A_27_367#_c_316_n N_VPWR_c_365_n 0.058048f $X=3.345 $Y=2.385 $X2=0
+ $Y2=0
cc_258 N_A_27_367#_c_318_n N_Y_M1004_s 0.00332344f $X=4.205 $Y=2.99 $X2=0 $Y2=0
cc_259 N_A_27_367#_M1008_d N_Y_c_438_n 0.00765997f $X=3.3 $Y=1.835 $X2=0 $Y2=0
cc_260 N_A_27_367#_c_316_n N_Y_c_438_n 0.0322441f $X=3.345 $Y=2.385 $X2=0 $Y2=0
cc_261 N_A_27_367#_c_348_p N_Y_c_438_n 0.0135577f $X=3.44 $Y=2.47 $X2=0 $Y2=0
cc_262 N_A_27_367#_c_318_n N_Y_c_444_n 0.0159805f $X=4.205 $Y=2.99 $X2=0 $Y2=0
cc_263 N_A_27_367#_c_297_n Y 0.0122795f $X=1.93 $Y=1.8 $X2=0 $Y2=0
cc_264 N_A_27_367#_c_316_n Y 0.0322159f $X=3.345 $Y=2.385 $X2=0 $Y2=0
cc_265 N_A_27_367#_c_295_n N_A_27_69#_c_502_n 0.00336159f $X=1.025 $Y=1.8 $X2=0
+ $Y2=0
cc_266 N_A_27_367#_c_297_n N_A_27_69#_c_509_n 0.00374355f $X=1.93 $Y=1.8 $X2=0
+ $Y2=0
cc_267 N_A_27_367#_c_297_n N_A_27_69#_c_498_n 0.0131402f $X=1.93 $Y=1.8 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_355_n N_Y_M1004_s 0.00225186f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_M1002_s N_Y_c_438_n 0.0087748f $X=2.35 $Y=1.835 $X2=0 $Y2=0
cc_270 N_VPWR_M1002_s Y 0.00337692f $X=2.35 $Y=1.835 $X2=0 $Y2=0
cc_271 N_VPWR_M1002_s Y 0.0068281f $X=2.35 $Y=1.835 $X2=0 $Y2=0
cc_272 N_Y_c_419_n N_A_27_69#_c_498_n 0.0370061f $X=2.5 $Y=0.69 $X2=0 $Y2=0
cc_273 N_Y_c_424_n N_A_27_69#_c_498_n 0.00981176f $X=2.562 $Y=1.17 $X2=0 $Y2=0
cc_274 N_Y_c_422_n N_VGND_M1006_d 0.00176461f $X=4.205 $Y=1.17 $X2=0 $Y2=0
cc_275 N_Y_c_421_n N_VGND_c_538_n 0.0228652f $X=3.44 $Y=0.49 $X2=0 $Y2=0
cc_276 N_Y_c_422_n N_VGND_c_538_n 0.0170777f $X=4.205 $Y=1.17 $X2=0 $Y2=0
cc_277 N_Y_c_423_n N_VGND_c_538_n 0.0229007f $X=4.3 $Y=0.49 $X2=0 $Y2=0
cc_278 N_Y_c_421_n N_VGND_c_539_n 0.00932149f $X=3.44 $Y=0.49 $X2=0 $Y2=0
cc_279 N_Y_c_423_n N_VGND_c_542_n 0.0127923f $X=4.3 $Y=0.49 $X2=0 $Y2=0
cc_280 N_Y_c_421_n N_VGND_c_543_n 0.00704609f $X=3.44 $Y=0.49 $X2=0 $Y2=0
cc_281 N_Y_c_423_n N_VGND_c_543_n 0.00966963f $X=4.3 $Y=0.49 $X2=0 $Y2=0
cc_282 N_Y_c_420_n N_A_282_69#_M1007_d 0.00256188f $X=3.345 $Y=1.17 $X2=0 $Y2=0
cc_283 N_Y_M1007_s N_A_282_69#_c_589_n 0.00271158f $X=2.375 $Y=0.345 $X2=0 $Y2=0
cc_284 N_Y_c_419_n N_A_282_69#_c_589_n 0.0214569f $X=2.5 $Y=0.69 $X2=0 $Y2=0
cc_285 N_Y_c_421_n N_A_282_69#_c_589_n 0.00536374f $X=3.44 $Y=0.49 $X2=0 $Y2=0
cc_286 N_Y_c_424_n N_A_282_69#_c_589_n 0.00286684f $X=2.562 $Y=1.17 $X2=0 $Y2=0
cc_287 N_Y_c_420_n N_A_282_69#_c_595_n 0.0213413f $X=3.345 $Y=1.17 $X2=0 $Y2=0
cc_288 N_A_27_69#_c_502_n N_VGND_M1009_d 0.00352133f $X=1.025 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_27_69#_c_496_n N_VGND_c_537_n 0.0134269f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_290 N_A_27_69#_c_502_n N_VGND_c_537_n 0.0170777f $X=1.025 $Y=0.955 $X2=0
+ $Y2=0
cc_291 N_A_27_69#_c_497_n N_VGND_c_537_n 0.0140502f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_292 N_A_27_69#_c_497_n N_VGND_c_539_n 0.0108528f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_293 N_A_27_69#_c_496_n N_VGND_c_541_n 0.0118048f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_294 N_A_27_69#_c_496_n N_VGND_c_543_n 0.00925234f $X=0.26 $Y=0.5 $X2=0 $Y2=0
cc_295 N_A_27_69#_c_497_n N_VGND_c_543_n 0.00850618f $X=1.12 $Y=0.5 $X2=0 $Y2=0
cc_296 N_A_27_69#_c_509_n N_A_282_69#_M1003_d 0.00333177f $X=1.815 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_297 N_A_27_69#_M1011_s N_A_282_69#_c_589_n 0.00263371f $X=1.84 $Y=0.345 $X2=0
+ $Y2=0
cc_298 N_A_27_69#_c_509_n N_A_282_69#_c_589_n 0.00396432f $X=1.815 $Y=0.955
+ $X2=0 $Y2=0
cc_299 N_A_27_69#_c_498_n N_A_282_69#_c_589_n 0.0205169f $X=1.98 $Y=0.7 $X2=0
+ $Y2=0
cc_300 N_A_27_69#_c_497_n N_A_282_69#_c_590_n 7.06642e-19 $X=1.12 $Y=0.5 $X2=0
+ $Y2=0
cc_301 N_A_27_69#_c_509_n N_A_282_69#_c_590_n 0.0130514f $X=1.815 $Y=0.955 $X2=0
+ $Y2=0
cc_302 N_VGND_c_538_n N_A_282_69#_c_589_n 0.00219498f $X=3.87 $Y=0.47 $X2=0
+ $Y2=0
cc_303 N_VGND_c_539_n N_A_282_69#_c_589_n 0.100214f $X=3.705 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_543_n N_A_282_69#_c_589_n 0.0565076f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_537_n N_A_282_69#_c_590_n 0.00244043f $X=0.69 $Y=0.575 $X2=0
+ $Y2=0
cc_306 N_VGND_c_539_n N_A_282_69#_c_590_n 0.0151402f $X=3.705 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_543_n N_A_282_69#_c_590_n 0.00838419f $X=4.56 $Y=0 $X2=0 $Y2=0
