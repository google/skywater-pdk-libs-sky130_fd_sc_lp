* File: sky130_fd_sc_lp__o221a_0.pxi.spice
* Created: Wed Sep  2 10:18:06 2020
* 
x_PM_SKY130_FD_SC_LP__O221A_0%C1 N_C1_M1005_g N_C1_M1008_g N_C1_c_82_n
+ N_C1_c_87_n C1 C1 C1 N_C1_c_84_n PM_SKY130_FD_SC_LP__O221A_0%C1
x_PM_SKY130_FD_SC_LP__O221A_0%B1 N_B1_M1007_g N_B1_c_125_n N_B1_M1003_g
+ N_B1_c_120_n N_B1_c_121_n N_B1_c_127_n B1 B1 N_B1_c_123_n N_B1_c_124_n
+ PM_SKY130_FD_SC_LP__O221A_0%B1
x_PM_SKY130_FD_SC_LP__O221A_0%B2 N_B2_c_166_n N_B2_M1000_g N_B2_M1002_g
+ N_B2_c_167_n N_B2_c_168_n N_B2_c_172_n N_B2_c_173_n B2 B2 N_B2_c_170_n
+ PM_SKY130_FD_SC_LP__O221A_0%B2
x_PM_SKY130_FD_SC_LP__O221A_0%A2 N_A2_M1011_g N_A2_c_218_n N_A2_M1001_g A2
+ N_A2_c_220_n PM_SKY130_FD_SC_LP__O221A_0%A2
x_PM_SKY130_FD_SC_LP__O221A_0%A1 N_A1_c_262_n N_A1_M1004_g N_A1_c_263_n
+ N_A1_M1009_g A1 A1 A1 N_A1_c_266_n PM_SKY130_FD_SC_LP__O221A_0%A1
x_PM_SKY130_FD_SC_LP__O221A_0%A_32_484# N_A_32_484#_M1008_s N_A_32_484#_M1005_s
+ N_A_32_484#_M1002_d N_A_32_484#_M1006_g N_A_32_484#_M1010_g
+ N_A_32_484#_c_310_n N_A_32_484#_c_315_n N_A_32_484#_c_316_n
+ N_A_32_484#_c_317_n N_A_32_484#_c_318_n N_A_32_484#_c_319_n
+ N_A_32_484#_c_311_n N_A_32_484#_c_320_n N_A_32_484#_c_321_n
+ N_A_32_484#_c_322_n PM_SKY130_FD_SC_LP__O221A_0%A_32_484#
x_PM_SKY130_FD_SC_LP__O221A_0%VPWR N_VPWR_M1005_d N_VPWR_M1004_d VPWR
+ N_VPWR_c_386_n N_VPWR_c_385_n N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_390_n
+ N_VPWR_c_391_n PM_SKY130_FD_SC_LP__O221A_0%VPWR
x_PM_SKY130_FD_SC_LP__O221A_0%X N_X_M1010_d N_X_M1006_d X X X X X X N_X_c_428_n
+ PM_SKY130_FD_SC_LP__O221A_0%X
x_PM_SKY130_FD_SC_LP__O221A_0%A_127_106# N_A_127_106#_M1008_d
+ N_A_127_106#_M1000_d N_A_127_106#_c_441_n N_A_127_106#_c_442_n
+ N_A_127_106#_c_443_n N_A_127_106#_c_444_n
+ PM_SKY130_FD_SC_LP__O221A_0%A_127_106#
x_PM_SKY130_FD_SC_LP__O221A_0%A_213_106# N_A_213_106#_M1007_d
+ N_A_213_106#_M1001_d N_A_213_106#_c_468_n N_A_213_106#_c_465_n
+ N_A_213_106#_c_466_n N_A_213_106#_c_467_n N_A_213_106#_c_493_n
+ PM_SKY130_FD_SC_LP__O221A_0%A_213_106#
x_PM_SKY130_FD_SC_LP__O221A_0%VGND N_VGND_M1001_s N_VGND_M1009_d N_VGND_c_507_n
+ N_VGND_c_508_n VGND N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n PM_SKY130_FD_SC_LP__O221A_0%VGND
cc_1 VNB N_C1_M1008_g 0.0441823f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_2 VNB N_C1_c_82_n 0.00272642f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.955
cc_3 VNB C1 0.0102582f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C1_c_84_n 0.0171195f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_5 VNB N_B1_c_120_n 0.0160695f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.12
cc_6 VNB N_B1_c_121_n 0.0109737f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB B1 0.0022502f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_8 VNB N_B1_c_123_n 0.0151833f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_9 VNB N_B1_c_124_n 0.0190955f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.295
cc_10 VNB N_B2_c_166_n 0.0174527f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.12
cc_11 VNB N_B2_c_167_n 0.0227996f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.12
cc_12 VNB N_B2_c_168_n 0.0169572f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_13 VNB B2 0.0036675f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_14 VNB N_B2_c_170_n 0.0136191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_M1011_g 0.0299127f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.74
cc_16 VNB N_A2_c_218_n 0.0198169f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.45
cc_17 VNB A2 0.0036257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_220_n 0.048424f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_19 VNB N_A1_c_262_n 0.0337813f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.12
cc_20 VNB N_A1_c_263_n 0.0235653f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_21 VNB N_A1_M1009_g 0.0228611f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_22 VNB A1 0.00984572f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_23 VNB N_A1_c_266_n 0.0176368f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_24 VNB N_A_32_484#_M1010_g 0.0698939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_32_484#_c_310_n 0.0358486f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_26 VNB N_A_32_484#_c_311_n 0.0152204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_385_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_28 VNB N_X_c_428_n 0.0703823f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_29 VNB N_A_127_106#_c_441_n 0.00185018f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_30 VNB N_A_127_106#_c_442_n 0.013022f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.955
cc_31 VNB N_A_127_106#_c_443_n 0.00850065f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.12
cc_32 VNB N_A_127_106#_c_444_n 0.00177055f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_33 VNB N_A_213_106#_c_465_n 0.0290778f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.955
cc_34 VNB N_A_213_106#_c_466_n 0.0025276f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.12
cc_35 VNB N_A_213_106#_c_467_n 0.00652135f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_36 VNB N_VGND_c_507_n 0.00918269f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.615
cc_37 VNB N_VGND_c_508_n 0.00506933f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_38 VNB N_VGND_c_509_n 0.0546731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_510_n 0.0179593f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.615
cc_40 VNB N_VGND_c_511_n 0.0175919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_512_n 0.233851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_513_n 0.0047828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_514_n 0.00632231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_C1_M1005_g 0.0331531f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.74
cc_45 VPB N_C1_c_82_n 0.0209026f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.955
cc_46 VPB N_C1_c_87_n 0.0166366f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.12
cc_47 VPB C1 0.00602346f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_48 VPB N_B1_c_125_n 0.0210949f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=0.74
cc_49 VPB N_B1_M1003_g 0.0236333f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.45
cc_50 VPB N_B1_c_127_n 0.021909f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_51 VPB B1 0.00149309f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_52 VPB N_B1_c_123_n 0.00644987f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.615
cc_53 VPB N_B2_M1002_g 0.0239748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B2_c_172_n 0.0187158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B2_c_173_n 0.0142742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB B2 0.0138709f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.615
cc_57 VPB N_B2_c_170_n 5.53722e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A2_M1011_g 0.0427043f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.74
cc_59 VPB N_A1_c_262_n 0.010697f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.12
cc_60 VPB N_A1_M1004_g 0.053257f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.74
cc_61 VPB A1 0.00597754f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_62 VPB N_A_32_484#_M1006_g 0.0241315f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.12
cc_63 VPB N_A_32_484#_M1010_g 0.0182628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_32_484#_c_310_n 0.0344056f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.615
cc_65 VPB N_A_32_484#_c_315_n 0.0217792f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.295
cc_66 VPB N_A_32_484#_c_316_n 0.0144294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_32_484#_c_317_n 0.00281149f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.035
cc_68 VPB N_A_32_484#_c_318_n 0.0124463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_32_484#_c_319_n 0.00434131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_32_484#_c_320_n 0.0107438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_32_484#_c_321_n 0.00265521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_32_484#_c_322_n 0.0525527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_386_n 0.017596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_385_n 0.0595996f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.615
cc_75 VPB N_VPWR_c_388_n 0.0163502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_389_n 0.0141708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_390_n 0.0372459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_391_n 0.0141708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.0147244f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.12
cc_80 VPB N_X_c_428_n 0.0510018f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.615
cc_81 N_C1_c_87_n N_B1_c_125_n 0.0116276f $X=0.55 $Y=2.12 $X2=0 $Y2=0
cc_82 N_C1_M1005_g N_B1_M1003_g 0.0105926f $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_83 N_C1_M1008_g N_B1_c_120_n 0.016786f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_84 C1 N_B1_c_121_n 6.39624e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_C1_M1005_g N_B1_c_127_n 0.00263136f $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_86 C1 B1 0.0542268f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_C1_c_84_n B1 4.97254e-19 $X=0.55 $Y=1.615 $X2=0 $Y2=0
cc_88 N_C1_c_82_n N_B1_c_123_n 0.0116276f $X=0.55 $Y=1.955 $X2=0 $Y2=0
cc_89 N_C1_M1008_g N_B1_c_124_n 0.00799155f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_90 C1 N_B1_c_124_n 0.0109583f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_91 N_C1_c_84_n N_B1_c_124_n 0.0116276f $X=0.55 $Y=1.615 $X2=0 $Y2=0
cc_92 N_C1_M1005_g N_A_32_484#_c_310_n 0.00798831f $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_93 N_C1_M1008_g N_A_32_484#_c_310_n 0.00925995f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_94 C1 N_A_32_484#_c_310_n 0.0843474f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_95 N_C1_c_84_n N_A_32_484#_c_310_n 0.0164925f $X=0.55 $Y=1.615 $X2=0 $Y2=0
cc_96 N_C1_M1005_g N_A_32_484#_c_315_n 3.34285e-19 $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_97 N_C1_M1005_g N_A_32_484#_c_316_n 0.0126866f $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_98 N_C1_c_87_n N_A_32_484#_c_316_n 0.0022467f $X=0.55 $Y=2.12 $X2=0 $Y2=0
cc_99 C1 N_A_32_484#_c_316_n 0.0327111f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_100 N_C1_c_84_n N_A_32_484#_c_311_n 0.00189998f $X=0.55 $Y=1.615 $X2=0 $Y2=0
cc_101 N_C1_M1005_g N_VPWR_c_385_n 0.00505747f $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_102 N_C1_M1005_g N_VPWR_c_388_n 0.00456975f $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_103 N_C1_M1005_g N_VPWR_c_389_n 0.0101427f $X=0.5 $Y=2.74 $X2=0 $Y2=0
cc_104 N_C1_M1008_g N_A_127_106#_c_441_n 0.00239908f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_105 C1 N_A_127_106#_c_441_n 0.0142149f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_106 N_C1_M1008_g N_A_127_106#_c_443_n 0.00133001f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_107 N_C1_M1008_g N_A_213_106#_c_468_n 0.0011612f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_108 C1 N_A_213_106#_c_468_n 0.00507389f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_109 C1 N_A_213_106#_c_466_n 0.0141177f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_110 N_C1_M1008_g N_VGND_c_509_n 0.00469064f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_111 N_C1_M1008_g N_VGND_c_512_n 0.0049649f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B1_c_120_n N_B2_c_166_n 0.0117709f $X=1.01 $Y=1.06 $X2=-0.19 $Y2=-0.245
cc_113 N_B1_M1003_g N_B2_M1002_g 0.0257062f $X=1.27 $Y=2.74 $X2=0 $Y2=0
cc_114 N_B1_c_121_n N_B2_c_167_n 0.00823713f $X=1.01 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B1_c_124_n N_B2_c_168_n 0.00872481f $X=1.15 $Y=1.545 $X2=0 $Y2=0
cc_116 N_B1_c_125_n N_B2_c_172_n 0.0257062f $X=1.15 $Y=2.02 $X2=0 $Y2=0
cc_117 N_B1_c_127_n N_B2_c_173_n 0.0257062f $X=1.15 $Y=2.215 $X2=0 $Y2=0
cc_118 B1 B2 0.0535915f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_119 N_B1_c_123_n B2 0.0042574f $X=1.12 $Y=1.71 $X2=0 $Y2=0
cc_120 B1 N_B2_c_170_n 8.14777e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_121 N_B1_c_123_n N_B2_c_170_n 0.0257062f $X=1.12 $Y=1.71 $X2=0 $Y2=0
cc_122 N_B1_M1003_g N_A_32_484#_c_316_n 0.0124863f $X=1.27 $Y=2.74 $X2=0 $Y2=0
cc_123 N_B1_c_127_n N_A_32_484#_c_316_n 0.00446867f $X=1.15 $Y=2.215 $X2=0 $Y2=0
cc_124 B1 N_A_32_484#_c_316_n 0.0236759f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_125 N_B1_M1003_g N_VPWR_c_385_n 0.00415982f $X=1.27 $Y=2.74 $X2=0 $Y2=0
cc_126 N_B1_M1003_g N_VPWR_c_389_n 0.0120228f $X=1.27 $Y=2.74 $X2=0 $Y2=0
cc_127 N_B1_M1003_g N_VPWR_c_390_n 0.00275188f $X=1.27 $Y=2.74 $X2=0 $Y2=0
cc_128 N_B1_c_120_n N_A_127_106#_c_441_n 0.00129069f $X=1.01 $Y=1.06 $X2=0 $Y2=0
cc_129 N_B1_c_120_n N_A_127_106#_c_442_n 0.0099303f $X=1.01 $Y=1.06 $X2=0 $Y2=0
cc_130 N_B1_c_120_n N_A_213_106#_c_468_n 0.00757357f $X=1.01 $Y=1.06 $X2=0 $Y2=0
cc_131 N_B1_c_121_n N_A_213_106#_c_468_n 0.00470114f $X=1.01 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_c_121_n N_A_213_106#_c_466_n 3.65144e-19 $X=1.01 $Y=1.21 $X2=0 $Y2=0
cc_133 B1 N_A_213_106#_c_466_n 0.0274232f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_134 N_B1_c_123_n N_A_213_106#_c_466_n 0.00206675f $X=1.12 $Y=1.71 $X2=0 $Y2=0
cc_135 N_B1_c_124_n N_A_213_106#_c_466_n 0.00550239f $X=1.15 $Y=1.545 $X2=0
+ $Y2=0
cc_136 N_B1_c_120_n N_VGND_c_509_n 6.5935e-19 $X=1.01 $Y=1.06 $X2=0 $Y2=0
cc_137 N_B2_M1002_g N_A2_M1011_g 0.0130199f $X=1.63 $Y=2.74 $X2=0 $Y2=0
cc_138 N_B2_c_167_n N_A2_M1011_g 0.0146353f $X=1.637 $Y=1.135 $X2=0 $Y2=0
cc_139 B2 N_A2_M1011_g 0.0237517f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_140 N_B2_c_170_n N_A2_M1011_g 0.0434316f $X=1.72 $Y=1.665 $X2=0 $Y2=0
cc_141 N_B2_c_166_n A2 0.00106002f $X=1.42 $Y=1.06 $X2=0 $Y2=0
cc_142 N_B2_c_166_n N_A2_c_220_n 0.00524924f $X=1.42 $Y=1.06 $X2=0 $Y2=0
cc_143 N_B2_c_167_n N_A2_c_220_n 0.0025227f $X=1.637 $Y=1.135 $X2=0 $Y2=0
cc_144 B2 N_A1_c_262_n 0.00394768f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_145 B2 A1 0.00699941f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_B2_M1002_g N_A_32_484#_c_316_n 0.00968356f $X=1.63 $Y=2.74 $X2=0 $Y2=0
cc_147 B2 N_A_32_484#_c_316_n 0.0163768f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 N_B2_M1002_g N_A_32_484#_c_317_n 2.11933e-19 $X=1.63 $Y=2.74 $X2=0 $Y2=0
cc_149 B2 N_A_32_484#_c_318_n 0.0138545f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_B2_c_173_n N_A_32_484#_c_321_n 0.00103873f $X=1.72 $Y=2.17 $X2=0 $Y2=0
cc_151 B2 N_A_32_484#_c_321_n 0.0308154f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_152 N_B2_M1002_g N_VPWR_c_385_n 0.00607506f $X=1.63 $Y=2.74 $X2=0 $Y2=0
cc_153 N_B2_M1002_g N_VPWR_c_389_n 0.0019633f $X=1.63 $Y=2.74 $X2=0 $Y2=0
cc_154 N_B2_M1002_g N_VPWR_c_390_n 0.00550375f $X=1.63 $Y=2.74 $X2=0 $Y2=0
cc_155 N_B2_c_166_n N_A_127_106#_c_442_n 0.0102969f $X=1.42 $Y=1.06 $X2=0 $Y2=0
cc_156 N_B2_c_167_n N_A_127_106#_c_442_n 9.65177e-19 $X=1.637 $Y=1.135 $X2=0
+ $Y2=0
cc_157 N_B2_c_166_n N_A_127_106#_c_444_n 0.00285484f $X=1.42 $Y=1.06 $X2=0 $Y2=0
cc_158 N_B2_c_167_n N_A_127_106#_c_444_n 0.005135f $X=1.637 $Y=1.135 $X2=0 $Y2=0
cc_159 N_B2_c_166_n N_A_213_106#_c_468_n 0.00778364f $X=1.42 $Y=1.06 $X2=0 $Y2=0
cc_160 N_B2_c_167_n N_A_213_106#_c_468_n 0.00669687f $X=1.637 $Y=1.135 $X2=0
+ $Y2=0
cc_161 N_B2_c_167_n N_A_213_106#_c_465_n 0.0132393f $X=1.637 $Y=1.135 $X2=0
+ $Y2=0
cc_162 N_B2_c_168_n N_A_213_106#_c_465_n 0.00940804f $X=1.72 $Y=1.5 $X2=0 $Y2=0
cc_163 B2 N_A_213_106#_c_465_n 0.0571803f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_B2_c_170_n N_A_213_106#_c_465_n 0.00446257f $X=1.72 $Y=1.665 $X2=0
+ $Y2=0
cc_165 N_B2_c_167_n N_A_213_106#_c_466_n 6.26939e-19 $X=1.637 $Y=1.135 $X2=0
+ $Y2=0
cc_166 N_B2_c_166_n N_VGND_c_507_n 4.89619e-19 $X=1.42 $Y=1.06 $X2=0 $Y2=0
cc_167 N_B2_c_166_n N_VGND_c_509_n 6.5935e-19 $X=1.42 $Y=1.06 $X2=0 $Y2=0
cc_168 N_A2_M1011_g N_A1_c_262_n 0.100838f $X=2.17 $Y=2.74 $X2=-0.19 $Y2=-0.245
cc_169 N_A2_c_220_n N_A1_c_262_n 3.86887e-19 $X=2.17 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A2_M1011_g N_A1_c_263_n 0.0107146f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_171 N_A2_c_218_n N_A1_M1009_g 0.0165387f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_172 N_A2_M1011_g A1 0.00106747f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_173 N_A2_c_220_n N_A1_c_266_n 0.00672429f $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_174 N_A2_M1011_g N_A_32_484#_c_317_n 2.11933e-19 $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_175 N_A2_M1011_g N_A_32_484#_c_318_n 0.00968356f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_176 N_A2_M1011_g N_VPWR_c_385_n 0.00607506f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_177 N_A2_M1011_g N_VPWR_c_390_n 0.00550375f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_178 N_A2_M1011_g N_VPWR_c_391_n 0.0019633f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_179 N_A2_c_218_n N_A_127_106#_c_444_n 0.00374581f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_180 A2 N_A_127_106#_c_444_n 0.0110882f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_181 N_A2_c_220_n N_A_127_106#_c_444_n 4.80875e-19 $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_182 A2 N_A_213_106#_c_468_n 0.00398688f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_183 N_A2_c_220_n N_A_213_106#_c_468_n 4.48906e-19 $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_184 N_A2_M1011_g N_A_213_106#_c_465_n 0.0114317f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_185 A2 N_A_213_106#_c_465_n 0.0261289f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_186 N_A2_c_220_n N_A_213_106#_c_465_n 0.0105531f $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_187 N_A2_M1011_g N_A_213_106#_c_467_n 0.00211994f $X=2.17 $Y=2.74 $X2=0 $Y2=0
cc_188 N_A2_c_218_n N_A_213_106#_c_467_n 0.0074121f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_189 A2 N_A_213_106#_c_467_n 0.018679f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_190 N_A2_c_220_n N_A_213_106#_c_467_n 0.00607792f $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_191 N_A2_c_218_n N_A_213_106#_c_493_n 0.00462441f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_192 N_A2_c_218_n N_VGND_c_507_n 0.00318258f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_193 A2 N_VGND_c_507_n 0.0189192f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_194 N_A2_c_220_n N_VGND_c_507_n 0.00634077f $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_195 N_A2_c_220_n N_VGND_c_509_n 0.00174653f $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_196 N_A2_c_218_n N_VGND_c_510_n 0.00533509f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_197 N_A2_c_220_n N_VGND_c_510_n 8.49756e-19 $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_198 N_A2_c_218_n N_VGND_c_512_n 0.0107754f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_199 A2 N_VGND_c_512_n 0.00508792f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_200 N_A2_c_220_n N_VGND_c_512_n 0.00354742f $X=2.17 $Y=0.93 $X2=0 $Y2=0
cc_201 N_A1_M1004_g N_A_32_484#_M1006_g 0.00796688f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_202 N_A1_c_262_n N_A_32_484#_M1010_g 0.00318036f $X=2.53 $Y=1.69 $X2=0 $Y2=0
cc_203 N_A1_M1004_g N_A_32_484#_M1010_g 0.00456308f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_204 N_A1_M1009_g N_A_32_484#_M1010_g 0.012159f $X=2.84 $Y=0.445 $X2=0 $Y2=0
cc_205 A1 N_A_32_484#_M1010_g 0.0084662f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_206 N_A1_c_266_n N_A_32_484#_M1010_g 0.0328666f $X=2.875 $Y=1.035 $X2=0 $Y2=0
cc_207 N_A1_c_262_n N_A_32_484#_c_318_n 0.00436128f $X=2.53 $Y=1.69 $X2=0 $Y2=0
cc_208 N_A1_M1004_g N_A_32_484#_c_318_n 0.0168902f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_209 A1 N_A_32_484#_c_318_n 0.00482528f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_210 N_A1_M1004_g N_A_32_484#_c_319_n 0.00471655f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_211 A1 N_A_32_484#_c_319_n 0.02783f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_212 N_A1_c_262_n N_A_32_484#_c_322_n 0.00305831f $X=2.53 $Y=1.69 $X2=0 $Y2=0
cc_213 N_A1_M1004_g N_A_32_484#_c_322_n 0.0126163f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_214 A1 N_A_32_484#_c_322_n 0.0022108f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_215 N_A1_M1004_g N_VPWR_c_385_n 0.00415982f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_216 N_A1_M1004_g N_VPWR_c_390_n 0.00275188f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_217 N_A1_M1004_g N_VPWR_c_391_n 0.0120228f $X=2.53 $Y=2.74 $X2=0 $Y2=0
cc_218 A1 N_X_c_428_n 0.082808f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_219 N_A1_c_262_n N_A_213_106#_c_465_n 0.00738962f $X=2.53 $Y=1.69 $X2=0 $Y2=0
cc_220 N_A1_c_263_n N_A_213_106#_c_465_n 0.00187592f $X=2.867 $Y=1.368 $X2=0
+ $Y2=0
cc_221 A1 N_A_213_106#_c_465_n 0.014702f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_222 N_A1_M1009_g N_A_213_106#_c_467_n 0.00403955f $X=2.84 $Y=0.445 $X2=0
+ $Y2=0
cc_223 A1 N_A_213_106#_c_467_n 0.031962f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_224 N_A1_c_266_n N_A_213_106#_c_467_n 0.00303913f $X=2.875 $Y=1.035 $X2=0
+ $Y2=0
cc_225 N_A1_c_266_n N_A_213_106#_c_493_n 0.00177447f $X=2.875 $Y=1.035 $X2=0
+ $Y2=0
cc_226 N_A1_M1009_g N_VGND_c_508_n 0.00190803f $X=2.84 $Y=0.445 $X2=0 $Y2=0
cc_227 A1 N_VGND_c_508_n 0.0257887f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_228 N_A1_c_266_n N_VGND_c_508_n 5.54583e-19 $X=2.875 $Y=1.035 $X2=0 $Y2=0
cc_229 N_A1_M1009_g N_VGND_c_510_n 0.00585385f $X=2.84 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A1_M1009_g N_VGND_c_512_n 0.00722301f $X=2.84 $Y=0.445 $X2=0 $Y2=0
cc_231 A1 N_VGND_c_512_n 0.00632984f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_232 N_A_32_484#_c_316_n N_VPWR_M1005_d 0.00721648f $X=1.735 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_233 N_A_32_484#_c_318_n N_VPWR_M1004_d 0.00700046f $X=2.935 $Y=2.47 $X2=0
+ $Y2=0
cc_234 N_A_32_484#_M1006_g N_VPWR_c_386_n 0.00456975f $X=3.3 $Y=2.74 $X2=0 $Y2=0
cc_235 N_A_32_484#_M1006_g N_VPWR_c_385_n 0.00846445f $X=3.3 $Y=2.74 $X2=0 $Y2=0
cc_236 N_A_32_484#_c_315_n N_VPWR_c_385_n 0.0102261f $X=0.285 $Y=2.565 $X2=0
+ $Y2=0
cc_237 N_A_32_484#_c_316_n N_VPWR_c_385_n 0.0244288f $X=1.735 $Y=2.47 $X2=0
+ $Y2=0
cc_238 N_A_32_484#_c_317_n N_VPWR_c_385_n 0.0127568f $X=1.9 $Y=2.56 $X2=0 $Y2=0
cc_239 N_A_32_484#_c_318_n N_VPWR_c_385_n 0.0197885f $X=2.935 $Y=2.47 $X2=0
+ $Y2=0
cc_240 N_A_32_484#_c_315_n N_VPWR_c_388_n 0.0188603f $X=0.285 $Y=2.565 $X2=0
+ $Y2=0
cc_241 N_A_32_484#_c_315_n N_VPWR_c_389_n 0.015234f $X=0.285 $Y=2.565 $X2=0
+ $Y2=0
cc_242 N_A_32_484#_c_316_n N_VPWR_c_389_n 0.0434634f $X=1.735 $Y=2.47 $X2=0
+ $Y2=0
cc_243 N_A_32_484#_c_317_n N_VPWR_c_389_n 0.00617689f $X=1.9 $Y=2.56 $X2=0 $Y2=0
cc_244 N_A_32_484#_c_317_n N_VPWR_c_390_n 0.0235393f $X=1.9 $Y=2.56 $X2=0 $Y2=0
cc_245 N_A_32_484#_M1006_g N_VPWR_c_391_n 0.0143164f $X=3.3 $Y=2.74 $X2=0 $Y2=0
cc_246 N_A_32_484#_c_317_n N_VPWR_c_391_n 0.00617689f $X=1.9 $Y=2.56 $X2=0 $Y2=0
cc_247 N_A_32_484#_c_318_n N_VPWR_c_391_n 0.0454171f $X=2.935 $Y=2.47 $X2=0
+ $Y2=0
cc_248 N_A_32_484#_c_322_n N_VPWR_c_391_n 0.00110425f $X=3.355 $Y=2.095 $X2=0
+ $Y2=0
cc_249 N_A_32_484#_c_316_n A_269_484# 0.00182165f $X=1.735 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_250 N_A_32_484#_c_318_n A_449_484# 0.00182165f $X=2.935 $Y=2.47 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_32_484#_M1006_g N_X_c_428_n 0.00906645f $X=3.3 $Y=2.74 $X2=0 $Y2=0
cc_252 N_A_32_484#_M1010_g N_X_c_428_n 0.0468213f $X=3.355 $Y=0.445 $X2=0 $Y2=0
cc_253 N_A_32_484#_c_318_n N_X_c_428_n 0.0140294f $X=2.935 $Y=2.47 $X2=0 $Y2=0
cc_254 N_A_32_484#_c_319_n N_X_c_428_n 0.0358398f $X=3.1 $Y=2.095 $X2=0 $Y2=0
cc_255 N_A_32_484#_M1010_g N_VGND_c_508_n 0.00335745f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_256 N_A_32_484#_c_311_n N_VGND_c_509_n 0.00724158f $X=0.345 $Y=0.74 $X2=0
+ $Y2=0
cc_257 N_A_32_484#_M1010_g N_VGND_c_511_n 0.00585385f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_258 N_A_32_484#_M1010_g N_VGND_c_512_n 0.0119989f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_259 N_A_32_484#_c_311_n N_VGND_c_512_n 0.0112095f $X=0.345 $Y=0.74 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_386_n X 0.0132849f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_c_385_n X 0.0121373f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_262 N_X_c_428_n N_VGND_c_511_n 0.0178245f $X=3.57 $Y=0.445 $X2=0 $Y2=0
cc_263 N_X_M1010_d N_VGND_c_512_n 0.00237743f $X=3.43 $Y=0.235 $X2=0 $Y2=0
cc_264 N_X_c_428_n N_VGND_c_512_n 0.012213f $X=3.57 $Y=0.445 $X2=0 $Y2=0
cc_265 N_A_127_106#_c_442_n N_A_213_106#_c_468_n 0.0207211f $X=1.54 $Y=0.347
+ $X2=0 $Y2=0
cc_266 N_A_127_106#_c_444_n N_A_213_106#_c_465_n 0.0100807f $X=1.635 $Y=0.74
+ $X2=0 $Y2=0
cc_267 N_A_127_106#_c_442_n N_VGND_c_507_n 0.0110576f $X=1.54 $Y=0.347 $X2=0
+ $Y2=0
cc_268 N_A_127_106#_c_444_n N_VGND_c_507_n 0.00827546f $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_269 N_A_127_106#_c_442_n N_VGND_c_509_n 0.0576428f $X=1.54 $Y=0.347 $X2=0
+ $Y2=0
cc_270 N_A_127_106#_c_443_n N_VGND_c_509_n 0.0157177f $X=0.87 $Y=0.347 $X2=0
+ $Y2=0
cc_271 N_A_127_106#_c_442_n N_VGND_c_512_n 0.0329941f $X=1.54 $Y=0.347 $X2=0
+ $Y2=0
cc_272 N_A_127_106#_c_443_n N_VGND_c_512_n 0.00854303f $X=0.87 $Y=0.347 $X2=0
+ $Y2=0
cc_273 N_A_213_106#_c_465_n N_VGND_c_507_n 2.78654e-19 $X=2.45 $Y=1.28 $X2=0
+ $Y2=0
cc_274 N_A_213_106#_c_493_n N_VGND_c_510_n 0.0149167f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_275 N_A_213_106#_M1001_d N_VGND_c_512_n 0.00226211f $X=2.485 $Y=0.235 $X2=0
+ $Y2=0
cc_276 N_A_213_106#_c_493_n N_VGND_c_512_n 0.0116779f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
