* File: sky130_fd_sc_lp__nor3b_4.pex.spice
* Created: Fri Aug 28 10:56:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3B_4%C_N 3 5 7 8 13
c28 3 0 5.52376e-20 $X=0.55 $Y=2.465
r29 11 13 3.31271 $w=2.91e-07 $l=2e-08 $layer=POLY_cond $X=0.53 $Y=1.35 $X2=0.55
+ $Y2=1.35
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.35 $X2=0.53 $Y2=1.35
r31 8 12 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.72 $Y=1.35 $X2=0.53
+ $Y2=1.35
r32 5 13 26.5017 $w=2.91e-07 $l=2.31571e-07 $layer=POLY_cond $X=0.71 $Y=1.185
+ $X2=0.55 $Y2=1.35
r33 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.71 $Y=1.185 $X2=0.71
+ $Y2=0.655
r34 1 13 18.2534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.515
+ $X2=0.55 $Y2=1.35
r35 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.55 $Y=1.515 $X2=0.55
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%A 1 3 6 8 10 13 15 17 20 22 24 27 31 32 34
+ 38 39 40
c90 39 0 5.52376e-20 $X=1.2 $Y=1.295
c91 32 0 2.20814e-20 $X=2.52 $Y=1.44
c92 27 0 1.73733e-19 $X=2.59 $Y=0.655
c93 20 0 6.17145e-20 $X=2.16 $Y=0.655
r94 55 56 12.2166 $w=4.34e-07 $l=1.1e-07 $layer=POLY_cond $X=2.16 $Y=1.5
+ $X2=2.27 $Y2=1.5
r95 51 53 16.659 $w=4.34e-07 $l=1.5e-07 $layer=POLY_cond $X=1.5 $Y=1.5 $X2=1.65
+ $Y2=1.5
r96 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.44 $X2=1.5 $Y2=1.44
r97 49 51 9.99539 $w=4.34e-07 $l=9e-08 $layer=POLY_cond $X=1.41 $Y=1.5 $X2=1.5
+ $Y2=1.5
r98 48 49 21.1014 $w=4.34e-07 $l=1.9e-07 $layer=POLY_cond $X=1.22 $Y=1.5
+ $X2=1.41 $Y2=1.5
r99 46 48 6.66359 $w=4.34e-07 $l=6e-08 $layer=POLY_cond $X=1.16 $Y=1.5 $X2=1.22
+ $Y2=1.5
r100 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.44 $X2=1.16 $Y2=1.44
r101 40 52 6.10117 $w=3.38e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.355
+ $X2=1.5 $Y2=1.355
r102 39 47 1.81413 $w=2.69e-07 $l=4e-08 $layer=LI1_cond $X=1.2 $Y=1.355 $X2=1.16
+ $Y2=1.355
r103 39 52 6.37438 $w=5.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.285 $Y=1.355
+ $X2=1.5 $Y2=1.355
r104 37 55 35.5392 $w=4.34e-07 $l=3.2e-07 $layer=POLY_cond $X=1.84 $Y=1.5
+ $X2=2.16 $Y2=1.5
r105 37 53 21.1014 $w=4.34e-07 $l=1.9e-07 $layer=POLY_cond $X=1.84 $Y=1.5
+ $X2=1.65 $Y2=1.5
r106 36 38 5.8358 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=1.84 $Y=1.355
+ $X2=1.955 $Y2=1.355
r107 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.84
+ $Y=1.44 $X2=1.84 $Y2=1.44
r108 34 40 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=1.355
+ $X2=1.68 $Y2=1.355
r109 34 36 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=1.785 $Y=1.355
+ $X2=1.84 $Y2=1.355
r110 32 58 7.77419 $w=4.34e-07 $l=7e-08 $layer=POLY_cond $X=2.52 $Y=1.5 $X2=2.59
+ $Y2=1.5
r111 32 56 27.765 $w=4.34e-07 $l=2.5e-07 $layer=POLY_cond $X=2.52 $Y=1.5
+ $X2=2.27 $Y2=1.5
r112 31 38 31.3318 $w=1.98e-07 $l=5.65e-07 $layer=LI1_cond $X=2.52 $Y=1.425
+ $X2=1.955 $Y2=1.425
r113 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.44 $X2=2.52 $Y2=1.44
r114 25 58 27.8684 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.59 $Y=1.275
+ $X2=2.59 $Y2=1.5
r115 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.59 $Y=1.275
+ $X2=2.59 $Y2=0.655
r116 22 56 27.8684 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.27 $Y=1.725
+ $X2=2.27 $Y2=1.5
r117 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.27 $Y=1.725
+ $X2=2.27 $Y2=2.465
r118 18 55 27.8684 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.16 $Y=1.275
+ $X2=2.16 $Y2=1.5
r119 18 20 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.16 $Y=1.275
+ $X2=2.16 $Y2=0.655
r120 15 37 27.8684 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.84 $Y=1.725
+ $X2=1.84 $Y2=1.5
r121 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.84 $Y=1.725
+ $X2=1.84 $Y2=2.465
r122 11 53 27.8684 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.65 $Y=1.275
+ $X2=1.65 $Y2=1.5
r123 11 13 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.65 $Y=1.275
+ $X2=1.65 $Y2=0.655
r124 8 49 27.8684 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.41 $Y=1.725
+ $X2=1.41 $Y2=1.5
r125 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.41 $Y=1.725
+ $X2=1.41 $Y2=2.465
r126 4 48 27.8684 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.22 $Y=1.275
+ $X2=1.22 $Y2=1.5
r127 4 6 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.22 $Y=1.275
+ $X2=1.22 $Y2=0.655
r128 1 46 19.9908 $w=4.34e-07 $l=3.01869e-07 $layer=POLY_cond $X=0.98 $Y=1.725
+ $X2=1.16 $Y2=1.5
r129 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.98 $Y=1.725
+ $X2=0.98 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%A_38_367# 1 2 9 11 13 16 18 20 23 25 27 30
+ 32 34 37 40 43 47 49 50 53 54 56 57
c135 30 0 6.17145e-20 $X=4.31 $Y=0.655
c136 23 0 1.73733e-19 $X=3.88 $Y=0.655
r137 67 68 24.6904 $w=4.49e-07 $l=2.3e-07 $layer=POLY_cond $X=4.08 $Y=1.49
+ $X2=4.31 $Y2=1.49
r138 66 67 21.4699 $w=4.49e-07 $l=2e-07 $layer=POLY_cond $X=3.88 $Y=1.49
+ $X2=4.08 $Y2=1.49
r139 65 66 24.6904 $w=4.49e-07 $l=2.3e-07 $layer=POLY_cond $X=3.65 $Y=1.49
+ $X2=3.88 $Y2=1.49
r140 64 65 21.4699 $w=4.49e-07 $l=2e-07 $layer=POLY_cond $X=3.45 $Y=1.49
+ $X2=3.65 $Y2=1.49
r141 63 64 24.6904 $w=4.49e-07 $l=2.3e-07 $layer=POLY_cond $X=3.22 $Y=1.49
+ $X2=3.45 $Y2=1.49
r142 60 63 17.1759 $w=4.49e-07 $l=1.6e-07 $layer=POLY_cond $X=3.06 $Y=1.49
+ $X2=3.22 $Y2=1.49
r143 60 61 4.29399 $w=4.49e-07 $l=4e-08 $layer=POLY_cond $X=3.06 $Y=1.49
+ $X2=3.02 $Y2=1.49
r144 59 60 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.06
+ $Y=1.42 $X2=3.06 $Y2=1.42
r145 54 70 9.66147 $w=4.49e-07 $l=9e-08 $layer=POLY_cond $X=4.42 $Y=1.49
+ $X2=4.51 $Y2=1.49
r146 54 68 11.8085 $w=4.49e-07 $l=1.1e-07 $layer=POLY_cond $X=4.42 $Y=1.49
+ $X2=4.31 $Y2=1.49
r147 53 54 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.42
+ $Y=1.42 $X2=4.42 $Y2=1.42
r148 51 59 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=1.415
+ $X2=2.98 $Y2=1.415
r149 51 53 83.4899 $w=1.78e-07 $l=1.355e-06 $layer=LI1_cond $X=3.065 $Y=1.415
+ $X2=4.42 $Y2=1.415
r150 49 59 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.98 $Y=1.505 $X2=2.98
+ $Y2=1.415
r151 49 50 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.98 $Y=1.505
+ $X2=2.98 $Y2=1.705
r152 48 57 2.79892 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.42 $Y=1.79
+ $X2=0.257 $Y2=1.79
r153 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.895 $Y=1.79
+ $X2=2.98 $Y2=1.705
r154 47 48 161.471 $w=1.68e-07 $l=2.475e-06 $layer=LI1_cond $X=2.895 $Y=1.79
+ $X2=0.42 $Y2=1.79
r155 43 45 32.9776 $w=3.23e-07 $l=9.3e-07 $layer=LI1_cond $X=0.257 $Y=1.98
+ $X2=0.257 $Y2=2.91
r156 41 57 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=1.875
+ $X2=0.257 $Y2=1.79
r157 41 43 3.72328 $w=3.23e-07 $l=1.05e-07 $layer=LI1_cond $X=0.257 $Y=1.875
+ $X2=0.257 $Y2=1.98
r158 40 57 3.67481 $w=2.52e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.185 $Y=1.705
+ $X2=0.257 $Y2=1.79
r159 40 56 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=0.185 $Y=1.705
+ $X2=0.185 $Y2=1.015
r160 35 56 10.9287 $w=4.83e-07 $l=2.42e-07 $layer=LI1_cond $X=0.337 $Y=0.773
+ $X2=0.337 $Y2=1.015
r161 35 37 8.70548 $w=4.83e-07 $l=3.53e-07 $layer=LI1_cond $X=0.337 $Y=0.773
+ $X2=0.337 $Y2=0.42
r162 32 70 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=4.51 $Y=1.725
+ $X2=4.51 $Y2=1.49
r163 32 34 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.51 $Y=1.725
+ $X2=4.51 $Y2=2.465
r164 28 68 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=4.31 $Y=1.255
+ $X2=4.31 $Y2=1.49
r165 28 30 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.31 $Y=1.255 $X2=4.31
+ $Y2=0.655
r166 25 67 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=4.08 $Y=1.725
+ $X2=4.08 $Y2=1.49
r167 25 27 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.08 $Y=1.725
+ $X2=4.08 $Y2=2.465
r168 21 66 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.88 $Y=1.255
+ $X2=3.88 $Y2=1.49
r169 21 23 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.88 $Y=1.255 $X2=3.88
+ $Y2=0.655
r170 18 65 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.65 $Y=1.725
+ $X2=3.65 $Y2=1.49
r171 18 20 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.65 $Y=1.725
+ $X2=3.65 $Y2=2.465
r172 14 64 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.45 $Y=1.255
+ $X2=3.45 $Y2=1.49
r173 14 16 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.45 $Y=1.255 $X2=3.45
+ $Y2=0.655
r174 11 63 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.22 $Y=1.725
+ $X2=3.22 $Y2=1.49
r175 11 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.22 $Y=1.725
+ $X2=3.22 $Y2=2.465
r176 7 61 28.7113 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.02 $Y=1.255
+ $X2=3.02 $Y2=1.49
r177 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.02 $Y=1.255 $X2=3.02
+ $Y2=0.655
r178 2 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.835 $X2=0.315 $Y2=2.91
r179 2 43 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.835 $X2=0.315 $Y2=1.98
r180 1 37 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.37
+ $Y=0.235 $X2=0.495 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%B 3 7 11 15 19 23 27 31 38 41 42 59 61 68 70
c86 27 0 1.73643e-19 $X=6.16 $Y=0.655
c87 15 0 6.04418e-20 $X=5.37 $Y=2.465
r88 61 68 0.117198 $w=2.93e-07 $l=3e-09 $layer=LI1_cond $X=5.523 $Y=1.357
+ $X2=5.52 $Y2=1.357
r89 58 59 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.16 $Y=1.42 $X2=6.23
+ $Y2=1.42
r90 55 56 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.73 $Y=1.42 $X2=5.8
+ $Y2=1.42
r91 52 53 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.3 $Y=1.42 $X2=5.37
+ $Y2=1.42
r92 50 52 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.03 $Y=1.42 $X2=5.3
+ $Y2=1.42
r93 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.03
+ $Y=1.42 $X2=5.03 $Y2=1.42
r94 48 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.94 $Y=1.42 $X2=5.03
+ $Y2=1.42
r95 46 48 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.87 $Y=1.42 $X2=4.94
+ $Y2=1.42
r96 42 70 6.19277 $w=2.93e-07 $l=1.06e-07 $layer=LI1_cond $X=5.564 $Y=1.357
+ $X2=5.67 $Y2=1.357
r97 42 61 1.6017 $w=2.93e-07 $l=4.1e-08 $layer=LI1_cond $X=5.564 $Y=1.357
+ $X2=5.523 $Y2=1.357
r98 42 68 1.6017 $w=2.93e-07 $l=4.1e-08 $layer=LI1_cond $X=5.479 $Y=1.357
+ $X2=5.52 $Y2=1.357
r99 41 42 17.1499 $w=2.93e-07 $l=4.39e-07 $layer=LI1_cond $X=5.04 $Y=1.357
+ $X2=5.479 $Y2=1.357
r100 41 51 0.390659 $w=2.93e-07 $l=1e-08 $layer=LI1_cond $X=5.04 $Y=1.357
+ $X2=5.03 $Y2=1.357
r101 39 58 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.05 $Y=1.42
+ $X2=6.16 $Y2=1.42
r102 39 56 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=6.05 $Y=1.42
+ $X2=5.8 $Y2=1.42
r103 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.05
+ $Y=1.42 $X2=6.05 $Y2=1.42
r104 36 55 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.71 $Y=1.42 $X2=5.73
+ $Y2=1.42
r105 36 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.71 $Y=1.42
+ $X2=5.37 $Y2=1.42
r106 35 38 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.71 $Y=1.42
+ $X2=6.05 $Y2=1.42
r107 35 70 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=5.71 $Y=1.42 $X2=5.67
+ $Y2=1.42
r108 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.71
+ $Y=1.42 $X2=5.71 $Y2=1.42
r109 29 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.585
+ $X2=6.23 $Y2=1.42
r110 29 31 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=6.23 $Y=1.585
+ $X2=6.23 $Y2=2.465
r111 25 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.255
+ $X2=6.16 $Y2=1.42
r112 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.16 $Y=1.255 $X2=6.16
+ $Y2=0.655
r113 21 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=1.585
+ $X2=5.8 $Y2=1.42
r114 21 23 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.8 $Y=1.585
+ $X2=5.8 $Y2=2.465
r115 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=1.255
+ $X2=5.73 $Y2=1.42
r116 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.73 $Y=1.255 $X2=5.73
+ $Y2=0.655
r117 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.37 $Y=1.585
+ $X2=5.37 $Y2=1.42
r118 13 15 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.37 $Y=1.585
+ $X2=5.37 $Y2=2.465
r119 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.3 $Y=1.255
+ $X2=5.3 $Y2=1.42
r120 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.3 $Y=1.255 $X2=5.3
+ $Y2=0.655
r121 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.94 $Y=1.585
+ $X2=4.94 $Y2=1.42
r122 5 7 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=4.94 $Y=1.585
+ $X2=4.94 $Y2=2.465
r123 1 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.87 $Y=1.255
+ $X2=4.87 $Y2=1.42
r124 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.87 $Y=1.255 $X2=4.87
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%VPWR 1 2 3 12 18 22 24 26 31 36 43 44 47 50
+ 53
r85 53 54 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r88 43 44 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=3.33
+ $X2=2.485 $Y2=3.33
r90 41 43 249.872 $w=1.68e-07 $l=3.83e-06 $layer=LI1_cond $X=2.65 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=3.33
+ $X2=1.625 $Y2=3.33
r95 37 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.79 $Y=3.33 $X2=2.16
+ $Y2=3.33
r96 36 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.485 $Y2=3.33
r97 36 39 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 35 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r101 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=3.33
+ $X2=0.765 $Y2=3.33
r102 32 34 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=3.33 $X2=1.2
+ $Y2=3.33
r103 31 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=3.33
+ $X2=1.625 $Y2=3.33
r104 31 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.46 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 29 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r107 26 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.765 $Y2=3.33
r108 26 28 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.24 $Y2=3.33
r109 24 44 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 24 54 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 20 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=3.245
+ $X2=2.485 $Y2=3.33
r112 20 22 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.485 $Y=3.245
+ $X2=2.485 $Y2=2.83
r113 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=3.245
+ $X2=1.625 $Y2=3.33
r114 16 18 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=1.625 $Y=3.245
+ $X2=1.625 $Y2=2.52
r115 12 15 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.765 $Y=2.19
+ $X2=0.765 $Y2=2.95
r116 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=3.245
+ $X2=0.765 $Y2=3.33
r117 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.765 $Y=3.245
+ $X2=0.765 $Y2=2.95
r118 3 22 600 $w=1.7e-07 $l=1.0627e-06 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=2.83
r119 2 18 300 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.52
r120 1 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.835 $X2=0.765 $Y2=2.95
r121 1 12 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.835 $X2=0.765 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%A_211_367# 1 2 3 4 13 15 17 21 23 25 31 38
+ 44
c65 23 0 6.04418e-20 $X=4.99 $Y=2.41
r66 40 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.155 $Y=2.115
+ $X2=5.155 $Y2=2.41
r67 38 40 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=5.155 $Y=2.11
+ $X2=5.155 $Y2=2.115
r68 35 36 4.62437 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=2.41
+ $X2=2.09 $Y2=2.495
r69 34 35 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=2.09 $Y=2.22 $X2=2.09
+ $Y2=2.41
r70 31 34 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=2.135
+ $X2=2.09 $Y2=2.22
r71 26 40 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=2.115
+ $X2=5.155 $Y2=2.115
r72 25 44 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.85 $Y=2.115
+ $X2=6.015 $Y2=2.115
r73 25 26 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=5.85 $Y=2.115
+ $X2=5.32 $Y2=2.115
r74 24 35 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.22 $Y=2.41 $X2=2.09
+ $Y2=2.41
r75 23 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=2.41
+ $X2=5.155 $Y2=2.41
r76 23 24 180.717 $w=1.68e-07 $l=2.77e-06 $layer=LI1_cond $X=4.99 $Y=2.41
+ $X2=2.22 $Y2=2.41
r77 21 36 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=2.055 $Y=2.56
+ $X2=2.055 $Y2=2.495
r78 18 30 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.29 $Y=2.135
+ $X2=1.195 $Y2=2.135
r79 17 31 2.89065 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=1.96 $Y=2.135
+ $X2=2.09 $Y2=2.135
r80 17 18 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=1.96 $Y=2.135
+ $X2=1.29 $Y2=2.135
r81 13 30 3.31928 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.195 $Y=2.225
+ $X2=1.195 $Y2=2.135
r82 13 15 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=1.195 $Y=2.225
+ $X2=1.195 $Y2=2.9
r83 4 44 300 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=2 $X=5.875
+ $Y=1.835 $X2=6.015 $Y2=2.11
r84 3 38 300 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=2 $X=5.015
+ $Y=1.835 $X2=5.155 $Y2=2.11
r85 2 34 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.22
r86 2 21 300 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=2 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.56
r87 1 30 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.835 $X2=1.195 $Y2=2.21
r88 1 15 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.835 $X2=1.195 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%A_576_367# 1 2 3 4 5 16 20 26 28 30 32 36 37
r47 35 36 7.66715 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=2.87
+ $X2=4.03 $Y2=2.87
r48 30 39 2.96959 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=6.48 $Y=2.885
+ $X2=6.48 $Y2=2.98
r49 30 32 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=6.48 $Y=2.885
+ $X2=6.48 $Y2=2.19
r50 29 37 5.05528 $w=1.95e-07 $l=9.74679e-08 $layer=LI1_cond $X=5.68 $Y=2.98
+ $X2=5.585 $Y2=2.975
r51 28 39 4.06365 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=6.35 $Y=2.98 $X2=6.48
+ $Y2=2.98
r52 28 29 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=6.35 $Y=2.98 $X2=5.68
+ $Y2=2.98
r53 24 37 1.43626 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=5.585 $Y=2.875
+ $X2=5.585 $Y2=2.975
r54 24 26 19.555 $w=1.88e-07 $l=3.35e-07 $layer=LI1_cond $X=5.585 $Y=2.875
+ $X2=5.585 $Y2=2.54
r55 23 36 38.5409 $w=1.98e-07 $l=6.95e-07 $layer=LI1_cond $X=4.725 $Y=2.975
+ $X2=4.03 $Y2=2.975
r56 20 37 5.05528 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=5.49 $Y=2.975
+ $X2=5.585 $Y2=2.975
r57 20 23 42.4227 $w=1.98e-07 $l=7.65e-07 $layer=LI1_cond $X=5.49 $Y=2.975
+ $X2=4.725 $Y2=2.975
r58 16 35 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=3.825 $Y=2.87
+ $X2=3.865 $Y2=2.87
r59 16 18 23.0489 $w=4.08e-07 $l=8.2e-07 $layer=LI1_cond $X=3.825 $Y=2.87
+ $X2=3.005 $Y2=2.87
r60 5 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.835 $X2=6.445 $Y2=2.91
r61 5 32 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.835 $X2=6.445 $Y2=2.19
r62 4 26 300 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_PDIFF $count=2 $X=5.445
+ $Y=1.835 $X2=5.585 $Y2=2.54
r63 3 23 600 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=1.835 $X2=4.725 $Y2=2.97
r64 2 35 600 $w=1.7e-07 $l=1.0627e-06 $layer=licon1_PDIFF $count=1 $X=3.725
+ $Y=1.835 $X2=3.865 $Y2=2.83
r65 1 18 600 $w=1.7e-07 $l=1.05565e-06 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.835 $X2=3.005 $Y2=2.83
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 41 43 49
+ 51 53 57 59 63 65 69 72 73 79 80 81 87
c132 81 0 1.73643e-19 $X=5.94 $Y=0.955
c133 73 0 1.73733e-19 $X=4.13 $Y=0.955
c134 69 0 1.73733e-19 $X=2.375 $Y=0.93
c135 43 0 2.20814e-20 $X=4.165 $Y=1.91
c136 41 0 6.17145e-20 $X=4 $Y=1.07
c137 35 0 6.17145e-20 $X=3.14 $Y=1.07
r138 86 87 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=6.51 $Y=1.675
+ $X2=6.51 $Y2=1.295
r139 85 87 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=6.51 $Y=1.155
+ $X2=6.51 $Y2=1.295
r140 81 83 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=5.94 $Y=0.955
+ $X2=5.94 $Y2=1.07
r141 81 82 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=0.955
+ $X2=5.94 $Y2=0.87
r142 78 79 7.41683 $w=4.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.295 $Y=1.91
+ $X2=4.4 $Y2=1.91
r143 73 75 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.13 $Y=0.955
+ $X2=4.13 $Y2=1.07
r144 73 74 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.955
+ $X2=4.13 $Y2=0.87
r145 69 70 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=2.34 $Y=0.93
+ $X2=2.34 $Y2=1.07
r146 68 69 3.94937 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.845
+ $X2=2.34 $Y2=0.93
r147 66 83 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.04 $Y=1.07 $X2=5.94
+ $Y2=1.07
r148 65 85 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.385 $Y=1.07
+ $X2=6.51 $Y2=1.155
r149 65 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.385 $Y=1.07
+ $X2=6.04 $Y2=1.07
r150 63 82 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=5.945 $Y=0.42
+ $X2=5.945 $Y2=0.87
r151 60 80 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.18 $Y=0.955
+ $X2=5.052 $Y2=0.955
r152 59 81 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.84 $Y=0.955 $X2=5.94
+ $Y2=0.955
r153 59 60 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.84 $Y=0.955
+ $X2=5.18 $Y2=0.955
r154 55 80 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.052 $Y=0.87
+ $X2=5.052 $Y2=0.955
r155 55 57 20.3372 $w=2.53e-07 $l=4.5e-07 $layer=LI1_cond $X=5.052 $Y=0.87
+ $X2=5.052 $Y2=0.42
r156 53 86 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=6.385 $Y=1.765
+ $X2=6.51 $Y2=1.675
r157 53 79 122.308 $w=1.78e-07 $l=1.985e-06 $layer=LI1_cond $X=6.385 $Y=1.765
+ $X2=4.4 $Y2=1.765
r158 52 73 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=0.955
+ $X2=4.13 $Y2=0.955
r159 51 80 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.925 $Y=0.955
+ $X2=5.052 $Y2=0.955
r160 51 52 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.925 $Y=0.955
+ $X2=4.26 $Y2=0.955
r161 49 74 20.3372 $w=2.53e-07 $l=4.5e-07 $layer=LI1_cond $X=4.127 $Y=0.42
+ $X2=4.127 $Y2=0.87
r162 43 78 3.3083 $w=4.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.165 $Y=1.91
+ $X2=4.295 $Y2=1.91
r163 43 45 18.5774 $w=4.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.165 $Y=1.91
+ $X2=3.435 $Y2=1.91
r164 42 72 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.33 $Y=1.07
+ $X2=3.235 $Y2=1.07
r165 41 75 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4 $Y=1.07 $X2=4.13
+ $Y2=1.07
r166 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4 $Y=1.07 $X2=3.33
+ $Y2=1.07
r167 37 72 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=0.985
+ $X2=3.235 $Y2=1.07
r168 37 39 32.9809 $w=1.88e-07 $l=5.65e-07 $layer=LI1_cond $X=3.235 $Y=0.985
+ $X2=3.235 $Y2=0.42
r169 36 70 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.47 $Y=1.07
+ $X2=2.34 $Y2=1.07
r170 35 72 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.14 $Y=1.07
+ $X2=3.235 $Y2=1.07
r171 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.14 $Y=1.07
+ $X2=2.47 $Y2=1.07
r172 33 68 21.2951 $w=2.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.355 $Y=0.42
+ $X2=2.355 $Y2=0.845
r173 29 69 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.21 $Y=0.93
+ $X2=2.34 $Y2=0.93
r174 29 30 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.21 $Y=0.93
+ $X2=1.57 $Y2=0.93
r175 25 30 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.437 $Y=0.845
+ $X2=1.57 $Y2=0.93
r176 25 27 18.4826 $w=2.63e-07 $l=4.25e-07 $layer=LI1_cond $X=1.437 $Y=0.845
+ $X2=1.437 $Y2=0.42
r177 8 78 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.155
+ $Y=1.835 $X2=4.295 $Y2=1.98
r178 7 45 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.835 $X2=3.435 $Y2=1.98
r179 6 63 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.805
+ $Y=0.235 $X2=5.945 $Y2=0.42
r180 5 57 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.945
+ $Y=0.235 $X2=5.085 $Y2=0.42
r181 4 49 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.955
+ $Y=0.235 $X2=4.095 $Y2=0.42
r182 3 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.095
+ $Y=0.235 $X2=3.235 $Y2=0.42
r183 2 69 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.235 $X2=2.375 $Y2=0.93
r184 2 33 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.235 $X2=2.375 $Y2=0.42
r185 1 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.295
+ $Y=0.235 $X2=1.435 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_4%VGND 1 2 3 4 5 6 7 24 28 30 34 38 42 46 48
+ 50 53 54 55 56 57 66 71 76 81 87 90 93 96 100
r105 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r106 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r107 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r108 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r109 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r110 85 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r111 85 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r112 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r113 82 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=5.515
+ $Y2=0
r114 82 84 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=6
+ $Y2=0
r115 81 99 4.60552 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=6.21 $Y=0 $X2=6.465
+ $Y2=0
r116 81 84 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.21 $Y=0 $X2=6
+ $Y2=0
r117 80 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r118 80 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r119 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r120 77 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.59
+ $Y2=0
r121 77 79 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=5.04 $Y2=0
r122 76 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.515
+ $Y2=0
r123 76 79 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.04
+ $Y2=0
r124 75 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r125 75 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r126 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r127 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.665
+ $Y2=0
r128 72 74 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.08
+ $Y2=0
r129 71 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.59
+ $Y2=0
r130 71 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.08
+ $Y2=0
r131 70 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r132 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r133 67 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.805
+ $Y2=0
r134 67 69 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=3.12
+ $Y2=0
r135 66 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.665
+ $Y2=0
r136 66 69 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.12
+ $Y2=0
r137 65 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r138 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r139 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r140 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r141 57 91 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r142 57 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r143 55 64 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.68
+ $Y2=0
r144 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.905
+ $Y2=0
r145 53 60 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.72
+ $Y2=0
r146 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.97
+ $Y2=0
r147 52 64 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=1.68 $Y2=0
r148 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.97
+ $Y2=0
r149 48 99 3.16065 $w=3.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.465 $Y2=0
r150 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0.38
r151 44 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0
r152 44 46 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0.56
r153 40 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0
r154 40 42 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0.56
r155 36 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=0.085
+ $X2=3.665 $Y2=0
r156 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.665 $Y=0.085
+ $X2=3.665 $Y2=0.36
r157 32 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=0.085
+ $X2=2.805 $Y2=0
r158 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.805 $Y=0.085
+ $X2=2.805 $Y2=0.36
r159 31 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.905
+ $Y2=0
r160 30 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.805
+ $Y2=0
r161 30 31 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.07
+ $Y2=0
r162 26 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=0.085
+ $X2=1.905 $Y2=0
r163 26 28 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.905 $Y=0.085
+ $X2=1.905 $Y2=0.545
r164 22 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0
r165 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0.38
r166 7 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.235
+ $Y=0.235 $X2=6.375 $Y2=0.38
r167 6 46 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=5.375
+ $Y=0.235 $X2=5.515 $Y2=0.56
r168 5 42 182 $w=1.7e-07 $l=4.1503e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.59 $Y2=0.56
r169 4 38 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.525
+ $Y=0.235 $X2=3.665 $Y2=0.36
r170 3 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.665
+ $Y=0.235 $X2=2.805 $Y2=0.36
r171 2 28 182 $w=1.7e-07 $l=3.89743e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.235 $X2=1.905 $Y2=0.545
r172 1 24 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=0.785
+ $Y=0.235 $X2=0.97 $Y2=0.38
.ends

