* File: sky130_fd_sc_lp__sdfxtp_4.pxi.spice
* Created: Fri Aug 28 11:30:57 2020
* 
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_91_123# N_A_91_123#_M1035_s N_A_91_123#_M1027_s
+ N_A_91_123#_M1037_g N_A_91_123#_M1007_g N_A_91_123#_c_245_n
+ N_A_91_123#_c_250_n N_A_91_123#_c_251_n N_A_91_123#_c_252_n
+ N_A_91_123#_c_246_n N_A_91_123#_c_247_n N_A_91_123#_c_248_n
+ PM_SKY130_FD_SC_LP__SDFXTP_4%A_91_123#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%D N_D_M1030_g N_D_M1020_g N_D_c_330_n N_D_c_331_n
+ N_D_c_332_n D D D D D N_D_c_334_n PM_SKY130_FD_SC_LP__SDFXTP_4%D
x_PM_SKY130_FD_SC_LP__SDFXTP_4%SCE N_SCE_c_382_n N_SCE_c_390_n N_SCE_c_391_n
+ N_SCE_M1035_g N_SCE_c_384_n N_SCE_c_385_n N_SCE_M1027_g N_SCE_c_393_n
+ N_SCE_M1016_g N_SCE_M1000_g N_SCE_c_395_n SCE SCE N_SCE_c_388_n
+ PM_SKY130_FD_SC_LP__SDFXTP_4%SCE
x_PM_SKY130_FD_SC_LP__SDFXTP_4%SCD N_SCD_M1001_g N_SCD_M1026_g SCD SCD
+ N_SCD_c_453_n PM_SKY130_FD_SC_LP__SDFXTP_4%SCD
x_PM_SKY130_FD_SC_LP__SDFXTP_4%CLK N_CLK_M1028_g N_CLK_M1031_g CLK CLK CLK
+ N_CLK_c_497_n PM_SKY130_FD_SC_LP__SDFXTP_4%CLK
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_641_123# N_A_641_123#_M1028_d
+ N_A_641_123#_M1031_d N_A_641_123#_M1006_g N_A_641_123#_c_540_n
+ N_A_641_123#_c_558_n N_A_641_123#_M1003_g N_A_641_123#_M1009_g
+ N_A_641_123#_M1022_g N_A_641_123#_M1023_g N_A_641_123#_M1034_g
+ N_A_641_123#_c_543_n N_A_641_123#_c_544_n N_A_641_123#_c_545_n
+ N_A_641_123#_c_561_n N_A_641_123#_c_546_n N_A_641_123#_c_547_n
+ N_A_641_123#_c_548_n N_A_641_123#_c_564_n N_A_641_123#_c_549_n
+ N_A_641_123#_c_550_n N_A_641_123#_c_630_p N_A_641_123#_c_566_n
+ N_A_641_123#_c_567_n N_A_641_123#_c_568_n N_A_641_123#_c_569_n
+ N_A_641_123#_c_570_n N_A_641_123#_c_571_n N_A_641_123#_c_551_n
+ N_A_641_123#_c_552_n N_A_641_123#_c_553_n N_A_641_123#_c_573_n
+ N_A_641_123#_c_554_n N_A_641_123#_c_574_n N_A_641_123#_c_555_n
+ N_A_641_123#_c_576_n N_A_641_123#_c_577_n N_A_641_123#_c_578_n
+ N_A_641_123#_c_556_n PM_SKY130_FD_SC_LP__SDFXTP_4%A_641_123#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_850_51# N_A_850_51#_M1006_d N_A_850_51#_M1003_d
+ N_A_850_51#_c_798_n N_A_850_51#_c_799_n N_A_850_51#_c_800_n
+ N_A_850_51#_c_801_n N_A_850_51#_M1008_g N_A_850_51#_c_780_n
+ N_A_850_51#_M1010_g N_A_850_51#_M1033_g N_A_850_51#_c_781_n
+ N_A_850_51#_c_782_n N_A_850_51#_c_783_n N_A_850_51#_M1032_g
+ N_A_850_51#_c_803_n N_A_850_51#_c_785_n N_A_850_51#_c_786_n
+ N_A_850_51#_c_787_n N_A_850_51#_c_788_n N_A_850_51#_c_789_n
+ N_A_850_51#_c_790_n N_A_850_51#_c_791_n N_A_850_51#_c_792_n
+ N_A_850_51#_c_793_n N_A_850_51#_c_794_n N_A_850_51#_c_795_n
+ N_A_850_51#_c_796_n N_A_850_51#_c_797_n PM_SKY130_FD_SC_LP__SDFXTP_4%A_850_51#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_1203_99# N_A_1203_99#_M1019_d
+ N_A_1203_99#_M1002_d N_A_1203_99#_c_955_n N_A_1203_99#_M1012_g
+ N_A_1203_99#_c_956_n N_A_1203_99#_c_957_n N_A_1203_99#_M1021_g
+ N_A_1203_99#_c_964_n N_A_1203_99#_c_958_n N_A_1203_99#_c_959_n
+ N_A_1203_99#_c_960_n N_A_1203_99#_c_961_n
+ PM_SKY130_FD_SC_LP__SDFXTP_4%A_1203_99#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_1053_125# N_A_1053_125#_M1009_d
+ N_A_1053_125#_M1008_d N_A_1053_125#_M1002_g N_A_1053_125#_c_1022_n
+ N_A_1053_125#_M1019_g N_A_1053_125#_c_1049_n N_A_1053_125#_c_1023_n
+ N_A_1053_125#_c_1024_n N_A_1053_125#_c_1028_n N_A_1053_125#_c_1025_n
+ N_A_1053_125#_c_1026_n PM_SKY130_FD_SC_LP__SDFXTP_4%A_1053_125#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_1673_409# N_A_1673_409#_M1013_d
+ N_A_1673_409#_M1015_d N_A_1673_409#_M1018_g N_A_1673_409#_M1029_g
+ N_A_1673_409#_c_1093_n N_A_1673_409#_M1005_g N_A_1673_409#_M1004_g
+ N_A_1673_409#_c_1095_n N_A_1673_409#_M1014_g N_A_1673_409#_M1011_g
+ N_A_1673_409#_c_1097_n N_A_1673_409#_M1017_g N_A_1673_409#_M1024_g
+ N_A_1673_409#_c_1099_n N_A_1673_409#_M1025_g N_A_1673_409#_M1036_g
+ N_A_1673_409#_c_1115_n N_A_1673_409#_c_1101_n N_A_1673_409#_c_1116_n
+ N_A_1673_409#_c_1102_n N_A_1673_409#_c_1103_n N_A_1673_409#_c_1104_n
+ N_A_1673_409#_c_1118_n N_A_1673_409#_c_1105_n N_A_1673_409#_c_1160_p
+ N_A_1673_409#_c_1106_n N_A_1673_409#_c_1107_n N_A_1673_409#_c_1120_n
+ N_A_1673_409#_c_1108_n PM_SKY130_FD_SC_LP__SDFXTP_4%A_1673_409#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_1475_449# N_A_1475_449#_M1033_d
+ N_A_1475_449#_M1023_d N_A_1475_449#_M1013_g N_A_1475_449#_M1015_g
+ N_A_1475_449#_c_1247_n N_A_1475_449#_c_1251_n N_A_1475_449#_c_1240_n
+ N_A_1475_449#_c_1241_n N_A_1475_449#_c_1242_n N_A_1475_449#_c_1233_n
+ N_A_1475_449#_c_1234_n N_A_1475_449#_c_1235_n N_A_1475_449#_c_1236_n
+ N_A_1475_449#_c_1237_n N_A_1475_449#_c_1238_n
+ PM_SKY130_FD_SC_LP__SDFXTP_4%A_1475_449#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%VPWR N_VPWR_M1027_d N_VPWR_M1001_d N_VPWR_M1003_s
+ N_VPWR_M1021_d N_VPWR_M1018_d N_VPWR_M1004_d N_VPWR_M1011_d N_VPWR_M1036_d
+ N_VPWR_c_1330_n N_VPWR_c_1331_n N_VPWR_c_1332_n N_VPWR_c_1333_n
+ N_VPWR_c_1334_n N_VPWR_c_1335_n N_VPWR_c_1336_n N_VPWR_c_1337_n
+ N_VPWR_c_1338_n N_VPWR_c_1339_n N_VPWR_c_1340_n N_VPWR_c_1341_n
+ N_VPWR_c_1342_n VPWR N_VPWR_c_1343_n N_VPWR_c_1344_n N_VPWR_c_1345_n
+ N_VPWR_c_1346_n N_VPWR_c_1347_n N_VPWR_c_1348_n N_VPWR_c_1349_n
+ N_VPWR_c_1350_n N_VPWR_c_1351_n N_VPWR_c_1329_n
+ PM_SKY130_FD_SC_LP__SDFXTP_4%VPWR
x_PM_SKY130_FD_SC_LP__SDFXTP_4%A_359_123# N_A_359_123#_M1030_d
+ N_A_359_123#_M1009_s N_A_359_123#_M1020_d N_A_359_123#_M1008_s
+ N_A_359_123#_c_1497_n N_A_359_123#_c_1508_n N_A_359_123#_c_1485_n
+ N_A_359_123#_c_1486_n N_A_359_123#_c_1500_n N_A_359_123#_c_1487_n
+ N_A_359_123#_c_1488_n N_A_359_123#_c_1491_n N_A_359_123#_c_1502_n
+ N_A_359_123#_c_1492_n N_A_359_123#_c_1493_n N_A_359_123#_c_1494_n
+ N_A_359_123#_c_1489_n PM_SKY130_FD_SC_LP__SDFXTP_4%A_359_123#
x_PM_SKY130_FD_SC_LP__SDFXTP_4%Q N_Q_M1005_s N_Q_M1017_s N_Q_M1004_s N_Q_M1024_s
+ N_Q_c_1604_n N_Q_c_1614_n N_Q_c_1605_n N_Q_c_1606_n N_Q_c_1611_n N_Q_c_1607_n
+ N_Q_c_1608_n N_Q_c_1644_n N_Q_c_1609_n N_Q_c_1613_n Q
+ PM_SKY130_FD_SC_LP__SDFXTP_4%Q
x_PM_SKY130_FD_SC_LP__SDFXTP_4%VGND N_VGND_M1035_d N_VGND_M1026_d N_VGND_M1006_s
+ N_VGND_M1012_d N_VGND_M1029_d N_VGND_M1005_d N_VGND_M1014_d N_VGND_M1025_d
+ N_VGND_c_1657_n N_VGND_c_1658_n N_VGND_c_1659_n N_VGND_c_1660_n
+ N_VGND_c_1661_n N_VGND_c_1662_n N_VGND_c_1663_n N_VGND_c_1664_n
+ N_VGND_c_1665_n N_VGND_c_1666_n N_VGND_c_1667_n N_VGND_c_1668_n
+ N_VGND_c_1669_n N_VGND_c_1670_n VGND N_VGND_c_1671_n N_VGND_c_1672_n
+ N_VGND_c_1673_n N_VGND_c_1674_n N_VGND_c_1675_n N_VGND_c_1676_n
+ N_VGND_c_1677_n N_VGND_c_1678_n N_VGND_c_1679_n N_VGND_c_1680_n
+ PM_SKY130_FD_SC_LP__SDFXTP_4%VGND
cc_1 VNB N_A_91_123#_M1037_g 0.0350636f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.825
cc_2 VNB N_A_91_123#_c_245_n 0.0338262f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.655
cc_3 VNB N_A_91_123#_c_246_n 0.0256617f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_4 VNB N_A_91_123#_c_247_n 0.0111876f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.74
cc_5 VNB N_A_91_123#_c_248_n 0.00643393f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.385
cc_6 VNB N_D_c_330_n 0.015223f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.825
cc_7 VNB N_D_c_331_n 0.028954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D_c_332_n 4.01051e-19 $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=2.295
cc_9 VNB D 0.00424774f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=2.775
cc_10 VNB N_D_c_334_n 0.021309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SCE_c_382_n 0.0114309f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.455
cc_12 VNB N_SCE_M1035_g 0.0357708f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.825
cc_13 VNB N_SCE_c_384_n 0.117423f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.825
cc_14 VNB N_SCE_c_385_n 0.0130655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_M1000_g 0.0358873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB SCE 0.00963678f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_17 VNB N_SCE_c_388_n 0.045125f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.385
cc_18 VNB N_SCD_M1026_g 0.0332046f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.575
cc_19 VNB SCD 0.00881234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_SCD_c_453_n 0.0243458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_CLK_M1028_g 0.0228383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB CLK 0.00803169f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=0.825
cc_23 VNB N_CLK_c_497_n 0.0458993f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.655
cc_24 VNB N_A_641_123#_c_540_n 0.00989061f $X=-0.19 $Y=-0.245 $X2=2.195
+ $Y2=2.295
cc_25 VNB N_A_641_123#_M1009_g 0.0384216f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.385
cc_26 VNB N_A_641_123#_M1034_g 0.0201337f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.74
cc_27 VNB N_A_641_123#_c_543_n 0.0245984f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.385
cc_28 VNB N_A_641_123#_c_544_n 0.0281355f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.78
cc_29 VNB N_A_641_123#_c_545_n 0.0157998f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.78
cc_30 VNB N_A_641_123#_c_546_n 0.00417537f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.295
cc_31 VNB N_A_641_123#_c_547_n 0.0322705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_641_123#_c_548_n 0.0133049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_641_123#_c_549_n 0.00519506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_641_123#_c_550_n 0.0105786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_641_123#_c_551_n 0.00232027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_641_123#_c_552_n 0.00656815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_641_123#_c_553_n 0.0336297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_641_123#_c_554_n 0.0195641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_641_123#_c_555_n 0.00125143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_641_123#_c_556_n 0.00699721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_850_51#_c_780_n 0.0142249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_850_51#_c_781_n 0.01501f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.13
cc_43 VNB N_A_850_51#_c_782_n 0.0200791f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.13
cc_44 VNB N_A_850_51#_c_783_n 0.0105409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_850_51#_M1032_g 0.00679484f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_46 VNB N_A_850_51#_c_785_n 0.00429032f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.385
cc_47 VNB N_A_850_51#_c_786_n 0.00173222f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.78
cc_48 VNB N_A_850_51#_c_787_n 0.0391846f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.74
cc_49 VNB N_A_850_51#_c_788_n 0.0322849f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.295
cc_50 VNB N_A_850_51#_c_789_n 0.0467218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_850_51#_c_790_n 0.00276968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_850_51#_c_791_n 0.00490135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_850_51#_c_792_n 0.00266181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_850_51#_c_793_n 0.0368157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_850_51#_c_794_n 0.00465208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_850_51#_c_795_n 0.0125204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_850_51#_c_796_n 0.0018547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_850_51#_c_797_n 0.0186885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1203_99#_c_955_n 0.0185607f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.575
cc_60 VNB N_A_1203_99#_c_956_n 0.0527279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1203_99#_c_957_n 0.00483516f $X=-0.19 $Y=-0.245 $X2=2.195
+ $Y2=2.295
cc_62 VNB N_A_1203_99#_c_958_n 0.00301506f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.385
cc_63 VNB N_A_1203_99#_c_959_n 0.00808115f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.13
cc_64 VNB N_A_1203_99#_c_960_n 0.0116464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1203_99#_c_961_n 0.00100926f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.74
cc_66 VNB N_A_1053_125#_M1002_g 0.0154527f $X=-0.19 $Y=-0.245 $X2=1.225
+ $Y2=0.825
cc_67 VNB N_A_1053_125#_c_1022_n 0.0228724f $X=-0.19 $Y=-0.245 $X2=2.195
+ $Y2=2.295
cc_68 VNB N_A_1053_125#_c_1023_n 0.0179924f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.13
cc_69 VNB N_A_1053_125#_c_1024_n 0.00248751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1053_125#_c_1025_n 0.00443666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1053_125#_c_1026_n 0.0408223f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.78
cc_72 VNB N_A_1673_409#_M1029_g 0.0556728f $X=-0.19 $Y=-0.245 $X2=2.195
+ $Y2=2.775
cc_73 VNB N_A_1673_409#_c_1093_n 0.0198708f $X=-0.19 $Y=-0.245 $X2=0.22
+ $Y2=0.965
cc_74 VNB N_A_1673_409#_M1004_g 0.00746195f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=2.13
cc_75 VNB N_A_1673_409#_c_1095_n 0.015823f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.13
cc_76 VNB N_A_1673_409#_M1011_g 0.00604603f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_77 VNB N_A_1673_409#_c_1097_n 0.0157986f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.74
cc_78 VNB N_A_1673_409#_M1024_g 0.00601356f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.78
cc_79 VNB N_A_1673_409#_c_1099_n 0.0186886f $X=-0.19 $Y=-0.245 $X2=1.225
+ $Y2=1.74
cc_80 VNB N_A_1673_409#_M1036_g 0.00684176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1673_409#_c_1101_n 0.00629726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1673_409#_c_1102_n 0.00523894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1673_409#_c_1103_n 5.05339e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1673_409#_c_1104_n 0.00413561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1673_409#_c_1105_n 0.0012629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1673_409#_c_1106_n 0.00210641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1673_409#_c_1107_n 0.0492998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1673_409#_c_1108_n 0.0749361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1475_449#_c_1233_n 0.00320151f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_90 VNB N_A_1475_449#_c_1234_n 0.00141535f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.74
cc_91 VNB N_A_1475_449#_c_1235_n 0.00739439f $X=-0.19 $Y=-0.245 $X2=0.7
+ $Y2=2.385
cc_92 VNB N_A_1475_449#_c_1236_n 0.0297096f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.78
cc_93 VNB N_A_1475_449#_c_1237_n 0.00250264f $X=-0.19 $Y=-0.245 $X2=1.105
+ $Y2=1.74
cc_94 VNB N_A_1475_449#_c_1238_n 0.0209327f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.13
cc_95 VNB N_VPWR_c_1329_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_359_123#_c_1485_n 0.0226651f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.13
cc_97 VNB N_A_359_123#_c_1486_n 0.00363574f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.13
cc_98 VNB N_A_359_123#_c_1487_n 0.00324f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_99 VNB N_A_359_123#_c_1488_n 0.00329631f $X=-0.19 $Y=-0.245 $X2=1.105
+ $Y2=1.74
cc_100 VNB N_A_359_123#_c_1489_n 0.00429971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_Q_c_1604_n 0.00120843f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=0.965
cc_102 VNB N_Q_c_1605_n 0.00309134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_Q_c_1606_n 0.00196569f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=0.8
cc_104 VNB N_Q_c_1607_n 0.00177567f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_105 VNB N_Q_c_1608_n 0.00120843f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.74
cc_106 VNB N_Q_c_1609_n 0.00834952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB Q 0.0270471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1657_n 0.00845358f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.8
cc_109 VNB N_VGND_c_1658_n 0.0185614f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.74
cc_110 VNB N_VGND_c_1659_n 0.015097f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.74
cc_111 VNB N_VGND_c_1660_n 0.00566471f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.295
cc_112 VNB N_VGND_c_1661_n 0.0150885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1662_n 6.48733e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1663_n 0.0108363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1664_n 0.024007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1665_n 0.0256963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1666_n 0.00463869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1667_n 0.0468185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1668_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1669_n 0.0177831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1670_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1671_n 0.0226891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1672_n 0.0497269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1673_n 0.0555935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1674_n 0.0150148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1675_n 0.0132031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1676_n 0.00526104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1677_n 0.0136387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1678_n 0.00494196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1679_n 0.00463869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1680_n 0.63247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VPB N_A_91_123#_M1007_g 0.0178384f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.775
cc_133 VPB N_A_91_123#_c_250_n 0.00970203f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=2.385
cc_134 VPB N_A_91_123#_c_251_n 0.00241045f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.13
cc_135 VPB N_A_91_123#_c_252_n 0.0366646f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.13
cc_136 VPB N_A_91_123#_c_247_n 0.0212111f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.74
cc_137 VPB N_A_91_123#_c_248_n 0.0792603f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.385
cc_138 VPB N_D_M1020_g 0.0471691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_D_c_332_n 0.0181608f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.295
cc_140 VPB D 0.00460875f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.775
cc_141 VPB N_SCE_c_382_n 0.0307597f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.455
cc_142 VPB N_SCE_c_390_n 0.0244481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_SCE_c_391_n 0.0109496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_SCE_M1027_g 0.0239857f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.775
cc_145 VPB N_SCE_c_393_n 0.0243446f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=0.965
cc_146 VPB N_SCE_M1016_g 0.0178524f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=2.3
cc_147 VPB N_SCE_c_395_n 0.00464609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_SCD_M1001_g 0.0526684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB SCD 0.0113022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_SCD_c_453_n 0.010611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_CLK_M1031_g 0.0467078f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=1.575
cc_152 VPB CLK 0.00944015f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=0.825
cc_153 VPB N_CLK_c_497_n 0.0278578f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.655
cc_154 VPB N_A_641_123#_c_540_n 0.0275806f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.295
cc_155 VPB N_A_641_123#_c_558_n 0.0236833f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.775
cc_156 VPB N_A_641_123#_M1022_g 0.0310773f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.13
cc_157 VPB N_A_641_123#_M1023_g 0.0231474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_641_123#_c_561_n 0.0259672f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.13
cc_159 VPB N_A_641_123#_c_546_n 0.0079092f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.295
cc_160 VPB N_A_641_123#_c_547_n 0.0347567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_641_123#_c_564_n 0.0120159f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_641_123#_c_550_n 0.0108059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_641_123#_c_566_n 0.0313594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_641_123#_c_567_n 0.00126212f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_641_123#_c_568_n 0.00313662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_641_123#_c_569_n 0.00445229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_641_123#_c_570_n 0.00288883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_641_123#_c_571_n 0.0138265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_641_123#_c_551_n 0.00583424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_641_123#_c_573_n 0.0107359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_641_123#_c_574_n 2.13598e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_641_123#_c_555_n 0.00129924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_641_123#_c_576_n 0.0115176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_641_123#_c_577_n 0.0445782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_641_123#_c_578_n 3.11147e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_850_51#_c_798_n 0.00823698f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=0.825
cc_177 VPB N_A_850_51#_c_799_n 0.0376076f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=0.825
cc_178 VPB N_A_850_51#_c_800_n 0.00963465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_850_51#_c_801_n 0.0215707f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.295
cc_180 VPB N_A_850_51#_M1032_g 0.0666802f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.8
cc_181 VPB N_A_850_51#_c_803_n 0.0163144f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.74
cc_182 VPB N_A_850_51#_c_786_n 0.0093955f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.78
cc_183 VPB N_A_850_51#_c_787_n 0.00558161f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.74
cc_184 VPB N_A_1203_99#_c_957_n 0.0159264f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.295
cc_185 VPB N_A_1203_99#_M1021_g 0.0196518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1203_99#_c_964_n 0.0182781f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.655
cc_187 VPB N_A_1203_99#_c_958_n 0.0106452f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=2.385
cc_188 VPB N_A_1203_99#_c_959_n 0.0010166f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.13
cc_189 VPB N_A_1053_125#_M1002_g 0.041205f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=0.825
cc_190 VPB N_A_1053_125#_c_1028_n 0.00237277f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.8
cc_191 VPB N_A_1053_125#_c_1025_n 0.00473481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_1673_409#_M1018_g 0.0221784f $X=-0.19 $Y=1.655 $X2=1.225
+ $Y2=0.825
cc_193 VPB N_A_1673_409#_M1029_g 0.0281423f $X=-0.19 $Y=1.655 $X2=2.195
+ $Y2=2.775
cc_194 VPB N_A_1673_409#_M1004_g 0.0243746f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=2.13
cc_195 VPB N_A_1673_409#_M1011_g 0.0181388f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.8
cc_196 VPB N_A_1673_409#_M1024_g 0.0181388f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.78
cc_197 VPB N_A_1673_409#_M1036_g 0.0227978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1673_409#_c_1115_n 0.00377318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_1673_409#_c_1116_n 0.00213052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1673_409#_c_1103_n 0.00460912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1673_409#_c_1118_n 0.0032847f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1673_409#_c_1107_n 0.00733038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1673_409#_c_1120_n 0.0413655f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1475_449#_M1015_g 0.0245437f $X=-0.19 $Y=1.655 $X2=2.195
+ $Y2=2.775
cc_205 VPB N_A_1475_449#_c_1240_n 0.0138498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1475_449#_c_1241_n 0.00864652f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=0.8
cc_207 VPB N_A_1475_449#_c_1242_n 0.00234017f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1475_449#_c_1234_n 3.97112e-19 $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.74
cc_209 VPB N_A_1475_449#_c_1236_n 0.00684763f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.78
cc_210 VPB N_VPWR_c_1330_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.8
cc_211 VPB N_VPWR_c_1331_n 0.00477979f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.74
cc_212 VPB N_VPWR_c_1332_n 0.0106013f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=1.74
cc_213 VPB N_VPWR_c_1333_n 0.0194722f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.295
cc_214 VPB N_VPWR_c_1334_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1335_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1336_n 0.0415885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1337_n 0.0391225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1338_n 0.00362538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1339_n 0.0186837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1340_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1341_n 0.0180085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1342_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1343_n 0.0284262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1344_n 0.0582658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1345_n 0.0471625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1346_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1347_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1348_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1349_n 0.0133114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1350_n 0.0223615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1351_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1329_n 0.100989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_359_123#_c_1487_n 0.00426002f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.8
cc_234 VPB N_A_359_123#_c_1491_n 0.0134144f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.78
cc_235 VPB N_A_359_123#_c_1492_n 0.00944765f $X=-0.19 $Y=1.655 $X2=2.215
+ $Y2=2.13
cc_236 VPB N_A_359_123#_c_1493_n 0.00182261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_359_123#_c_1494_n 0.00282953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_359_123#_c_1489_n 0.00530232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_Q_c_1611_n 0.00834361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_Q_c_1607_n 0.00408124f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.8
cc_241 VPB N_Q_c_1613_n 0.0136311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 N_A_91_123#_M1007_g N_D_M1020_g 0.0258655f $X=2.195 $Y=2.775 $X2=0 $Y2=0
cc_243 N_A_91_123#_c_250_n N_D_M1020_g 0.013302f $X=2.05 $Y=2.385 $X2=0 $Y2=0
cc_244 N_A_91_123#_c_251_n N_D_M1020_g 0.0017201f $X=2.215 $Y=2.13 $X2=0 $Y2=0
cc_245 N_A_91_123#_c_252_n N_D_M1020_g 0.0202023f $X=2.215 $Y=2.13 $X2=0 $Y2=0
cc_246 N_A_91_123#_c_247_n N_D_M1020_g 0.00230676f $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_247 N_A_91_123#_c_248_n N_D_M1020_g 0.00178503f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_248 N_A_91_123#_M1037_g N_D_c_330_n 0.0202689f $X=1.225 $Y=0.825 $X2=0 $Y2=0
cc_249 N_A_91_123#_c_247_n N_D_c_331_n 0.0183158f $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_250 N_A_91_123#_c_250_n N_D_c_332_n 6.29193e-19 $X=2.05 $Y=2.385 $X2=0 $Y2=0
cc_251 N_A_91_123#_c_247_n N_D_c_332_n 0.0048037f $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_252 N_A_91_123#_c_248_n N_D_c_332_n 5.6331e-19 $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_253 N_A_91_123#_M1037_g D 0.00949373f $X=1.225 $Y=0.825 $X2=0 $Y2=0
cc_254 N_A_91_123#_c_250_n D 0.021517f $X=2.05 $Y=2.385 $X2=0 $Y2=0
cc_255 N_A_91_123#_c_251_n D 0.00814041f $X=2.215 $Y=2.13 $X2=0 $Y2=0
cc_256 N_A_91_123#_c_252_n D 5.22061e-19 $X=2.215 $Y=2.13 $X2=0 $Y2=0
cc_257 N_A_91_123#_c_247_n D 4.70389e-19 $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_258 N_A_91_123#_c_248_n D 0.0305764f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_259 N_A_91_123#_M1037_g N_D_c_334_n 0.0183158f $X=1.225 $Y=0.825 $X2=0 $Y2=0
cc_260 N_A_91_123#_M1037_g N_SCE_c_382_n 0.00249596f $X=1.225 $Y=0.825 $X2=0
+ $Y2=0
cc_261 N_A_91_123#_c_247_n N_SCE_c_382_n 0.010041f $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_262 N_A_91_123#_c_248_n N_SCE_c_382_n 0.0292512f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_263 N_A_91_123#_c_248_n N_SCE_c_390_n 0.0199549f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_264 N_A_91_123#_c_248_n N_SCE_c_391_n 0.00862116f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_265 N_A_91_123#_M1037_g N_SCE_M1035_g 0.0192593f $X=1.225 $Y=0.825 $X2=0
+ $Y2=0
cc_266 N_A_91_123#_c_245_n N_SCE_M1035_g 0.00430998f $X=0.22 $Y=1.655 $X2=0
+ $Y2=0
cc_267 N_A_91_123#_M1037_g N_SCE_c_384_n 0.0103421f $X=1.225 $Y=0.825 $X2=0
+ $Y2=0
cc_268 N_A_91_123#_c_248_n N_SCE_M1027_g 0.0140918f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_269 N_A_91_123#_c_247_n N_SCE_c_393_n 0.001091f $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_270 N_A_91_123#_c_248_n N_SCE_c_393_n 0.00955477f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_271 N_A_91_123#_c_250_n N_SCE_M1016_g 0.0151157f $X=2.05 $Y=2.385 $X2=0 $Y2=0
cc_272 N_A_91_123#_c_248_n N_SCE_M1016_g 0.00109656f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_273 N_A_91_123#_c_247_n N_SCE_c_395_n 0.0214451f $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_274 N_A_91_123#_c_248_n N_SCE_c_395_n 0.0040142f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_275 N_A_91_123#_M1037_g SCE 0.0184551f $X=1.225 $Y=0.825 $X2=0 $Y2=0
cc_276 N_A_91_123#_c_245_n SCE 0.0263181f $X=0.22 $Y=1.655 $X2=0 $Y2=0
cc_277 N_A_91_123#_c_246_n SCE 0.0140226f $X=0.58 $Y=0.8 $X2=0 $Y2=0
cc_278 N_A_91_123#_c_247_n SCE 0.00523191f $X=1.105 $Y=1.74 $X2=0 $Y2=0
cc_279 N_A_91_123#_c_248_n SCE 0.0637348f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_280 N_A_91_123#_M1037_g N_SCE_c_388_n 0.00465083f $X=1.225 $Y=0.825 $X2=0
+ $Y2=0
cc_281 N_A_91_123#_c_245_n N_SCE_c_388_n 0.0151819f $X=0.22 $Y=1.655 $X2=0 $Y2=0
cc_282 N_A_91_123#_c_246_n N_SCE_c_388_n 0.00816907f $X=0.58 $Y=0.8 $X2=0 $Y2=0
cc_283 N_A_91_123#_c_248_n N_SCE_c_388_n 0.00272112f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_284 N_A_91_123#_M1007_g N_SCD_M1001_g 0.0356704f $X=2.195 $Y=2.775 $X2=0
+ $Y2=0
cc_285 N_A_91_123#_c_250_n N_SCD_M1001_g 5.02752e-19 $X=2.05 $Y=2.385 $X2=0
+ $Y2=0
cc_286 N_A_91_123#_c_251_n N_SCD_M1001_g 7.69607e-19 $X=2.215 $Y=2.13 $X2=0
+ $Y2=0
cc_287 N_A_91_123#_c_252_n N_SCD_M1001_g 0.0203469f $X=2.215 $Y=2.13 $X2=0 $Y2=0
cc_288 N_A_91_123#_c_250_n SCD 0.00396215f $X=2.05 $Y=2.385 $X2=0 $Y2=0
cc_289 N_A_91_123#_c_251_n SCD 0.0214873f $X=2.215 $Y=2.13 $X2=0 $Y2=0
cc_290 N_A_91_123#_c_252_n SCD 0.00486195f $X=2.215 $Y=2.13 $X2=0 $Y2=0
cc_291 N_A_91_123#_c_248_n N_VPWR_M1027_d 0.00178184f $X=0.7 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_91_123#_c_250_n N_VPWR_c_1330_n 0.00188374f $X=2.05 $Y=2.385 $X2=0
+ $Y2=0
cc_293 N_A_91_123#_c_248_n N_VPWR_c_1330_n 0.0163125f $X=0.7 $Y=2.385 $X2=0
+ $Y2=0
cc_294 N_A_91_123#_M1007_g N_VPWR_c_1337_n 0.0037886f $X=2.195 $Y=2.775 $X2=0
+ $Y2=0
cc_295 N_A_91_123#_c_248_n N_VPWR_c_1343_n 0.027891f $X=0.7 $Y=2.385 $X2=0 $Y2=0
cc_296 N_A_91_123#_M1027_s N_VPWR_c_1329_n 0.0025987f $X=0.635 $Y=2.455 $X2=0
+ $Y2=0
cc_297 N_A_91_123#_M1007_g N_VPWR_c_1329_n 0.00564534f $X=2.195 $Y=2.775 $X2=0
+ $Y2=0
cc_298 N_A_91_123#_c_250_n N_VPWR_c_1329_n 0.0144288f $X=2.05 $Y=2.385 $X2=0
+ $Y2=0
cc_299 N_A_91_123#_c_248_n N_VPWR_c_1329_n 0.0327174f $X=0.7 $Y=2.385 $X2=0
+ $Y2=0
cc_300 N_A_91_123#_c_250_n A_296_491# 0.00196273f $X=2.05 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_301 N_A_91_123#_c_250_n N_A_359_123#_M1020_d 0.00173028f $X=2.05 $Y=2.385
+ $X2=0 $Y2=0
cc_302 N_A_91_123#_M1007_g N_A_359_123#_c_1497_n 0.0129223f $X=2.195 $Y=2.775
+ $X2=0 $Y2=0
cc_303 N_A_91_123#_c_250_n N_A_359_123#_c_1497_n 0.025551f $X=2.05 $Y=2.385
+ $X2=0 $Y2=0
cc_304 N_A_91_123#_c_252_n N_A_359_123#_c_1497_n 0.00231433f $X=2.215 $Y=2.13
+ $X2=0 $Y2=0
cc_305 N_A_91_123#_M1007_g N_A_359_123#_c_1500_n 0.00298028f $X=2.195 $Y=2.775
+ $X2=0 $Y2=0
cc_306 N_A_91_123#_c_251_n N_A_359_123#_c_1487_n 0.00537829f $X=2.215 $Y=2.13
+ $X2=0 $Y2=0
cc_307 N_A_91_123#_c_250_n N_A_359_123#_c_1502_n 0.00134746f $X=2.05 $Y=2.385
+ $X2=0 $Y2=0
cc_308 N_A_91_123#_M1007_g N_A_359_123#_c_1492_n 0.00112861f $X=2.195 $Y=2.775
+ $X2=0 $Y2=0
cc_309 N_A_91_123#_c_250_n N_A_359_123#_c_1492_n 0.0135841f $X=2.05 $Y=2.385
+ $X2=0 $Y2=0
cc_310 N_A_91_123#_c_251_n N_A_359_123#_c_1492_n 0.0118139f $X=2.215 $Y=2.13
+ $X2=0 $Y2=0
cc_311 N_A_91_123#_c_252_n N_A_359_123#_c_1492_n 9.68269e-19 $X=2.215 $Y=2.13
+ $X2=0 $Y2=0
cc_312 N_A_91_123#_M1037_g N_VGND_c_1657_n 0.00911227f $X=1.225 $Y=0.825 $X2=0
+ $Y2=0
cc_313 N_A_91_123#_c_245_n N_VGND_c_1657_n 3.17897e-19 $X=0.22 $Y=1.655 $X2=0
+ $Y2=0
cc_314 N_A_91_123#_c_246_n N_VGND_c_1665_n 0.0101333f $X=0.58 $Y=0.8 $X2=0 $Y2=0
cc_315 N_A_91_123#_M1037_g N_VGND_c_1680_n 7.6887e-19 $X=1.225 $Y=0.825 $X2=0
+ $Y2=0
cc_316 N_A_91_123#_c_246_n N_VGND_c_1680_n 0.0159967f $X=0.58 $Y=0.8 $X2=0 $Y2=0
cc_317 N_D_c_330_n N_SCE_c_384_n 0.0091524f $X=1.675 $Y=1.145 $X2=0 $Y2=0
cc_318 D N_SCE_c_384_n 0.00411261f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_319 N_D_M1020_g N_SCE_c_393_n 0.0697571f $X=1.765 $Y=2.775 $X2=0 $Y2=0
cc_320 N_D_c_330_n N_SCE_M1000_g 0.0133867f $X=1.675 $Y=1.145 $X2=0 $Y2=0
cc_321 D N_SCE_M1000_g 0.00182937f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_322 N_D_c_334_n N_SCE_M1000_g 4.64914e-19 $X=1.675 $Y=1.31 $X2=0 $Y2=0
cc_323 D SCE 0.0272161f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_324 N_D_c_334_n SCE 0.0020084f $X=1.675 $Y=1.31 $X2=0 $Y2=0
cc_325 N_D_c_331_n SCD 0.00572464f $X=1.675 $Y=1.65 $X2=0 $Y2=0
cc_326 D SCD 0.0330292f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_327 N_D_c_331_n N_SCD_c_453_n 0.00419322f $X=1.675 $Y=1.65 $X2=0 $Y2=0
cc_328 D N_SCD_c_453_n 2.04755e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_329 N_D_M1020_g N_VPWR_c_1330_n 0.00266076f $X=1.765 $Y=2.775 $X2=0 $Y2=0
cc_330 N_D_M1020_g N_VPWR_c_1337_n 0.00550964f $X=1.765 $Y=2.775 $X2=0 $Y2=0
cc_331 N_D_M1020_g N_VPWR_c_1329_n 0.00626038f $X=1.765 $Y=2.775 $X2=0 $Y2=0
cc_332 N_D_M1020_g N_A_359_123#_c_1497_n 0.00589211f $X=1.765 $Y=2.775 $X2=0
+ $Y2=0
cc_333 N_D_c_330_n N_A_359_123#_c_1508_n 0.00248287f $X=1.675 $Y=1.145 $X2=0
+ $Y2=0
cc_334 D N_A_359_123#_c_1508_n 0.0234018f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_335 N_D_c_330_n N_A_359_123#_c_1486_n 8.55115e-19 $X=1.675 $Y=1.145 $X2=0
+ $Y2=0
cc_336 D N_A_359_123#_c_1486_n 0.0140876f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_337 N_D_c_334_n N_A_359_123#_c_1486_n 0.00146044f $X=1.675 $Y=1.31 $X2=0
+ $Y2=0
cc_338 N_D_c_330_n N_VGND_c_1657_n 4.45665e-19 $X=1.675 $Y=1.145 $X2=0 $Y2=0
cc_339 D N_VGND_c_1657_n 0.023196f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_340 D N_VGND_c_1667_n 0.00787289f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_341 D N_VGND_c_1680_n 0.00793227f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_342 D A_260_123# 0.00485688f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_343 N_SCE_M1000_g N_SCD_M1026_g 0.0418196f $X=2.34 $Y=0.825 $X2=0 $Y2=0
cc_344 N_SCE_M1000_g SCD 9.71168e-19 $X=2.34 $Y=0.825 $X2=0 $Y2=0
cc_345 N_SCE_M1027_g N_VPWR_c_1330_n 0.0157896f $X=0.975 $Y=2.775 $X2=0 $Y2=0
cc_346 N_SCE_c_393_n N_VPWR_c_1330_n 4.99926e-19 $X=1.33 $Y=2.19 $X2=0 $Y2=0
cc_347 N_SCE_M1016_g N_VPWR_c_1330_n 0.0137053f $X=1.405 $Y=2.775 $X2=0 $Y2=0
cc_348 N_SCE_M1016_g N_VPWR_c_1337_n 0.00486043f $X=1.405 $Y=2.775 $X2=0 $Y2=0
cc_349 N_SCE_M1027_g N_VPWR_c_1343_n 0.00486043f $X=0.975 $Y=2.775 $X2=0 $Y2=0
cc_350 N_SCE_M1027_g N_VPWR_c_1329_n 0.00605869f $X=0.975 $Y=2.775 $X2=0 $Y2=0
cc_351 N_SCE_M1016_g N_VPWR_c_1329_n 0.00449316f $X=1.405 $Y=2.775 $X2=0 $Y2=0
cc_352 N_SCE_M1016_g N_A_359_123#_c_1497_n 8.88788e-19 $X=1.405 $Y=2.775 $X2=0
+ $Y2=0
cc_353 N_SCE_c_384_n N_A_359_123#_c_1508_n 0.0033819f $X=2.265 $Y=0.2 $X2=0
+ $Y2=0
cc_354 N_SCE_M1000_g N_A_359_123#_c_1508_n 0.00604792f $X=2.34 $Y=0.825 $X2=0
+ $Y2=0
cc_355 N_SCE_M1000_g N_A_359_123#_c_1485_n 0.013329f $X=2.34 $Y=0.825 $X2=0
+ $Y2=0
cc_356 N_SCE_M1035_g N_VGND_c_1657_n 0.0255639f $X=0.795 $Y=0.825 $X2=0 $Y2=0
cc_357 N_SCE_c_384_n N_VGND_c_1657_n 0.01895f $X=2.265 $Y=0.2 $X2=0 $Y2=0
cc_358 N_SCE_c_385_n N_VGND_c_1657_n 0.00433435f $X=0.87 $Y=0.2 $X2=0 $Y2=0
cc_359 SCE N_VGND_c_1657_n 0.0229042f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_360 N_SCE_c_384_n N_VGND_c_1658_n 0.0104303f $X=2.265 $Y=0.2 $X2=0 $Y2=0
cc_361 N_SCE_M1000_g N_VGND_c_1658_n 0.00164631f $X=2.34 $Y=0.825 $X2=0 $Y2=0
cc_362 N_SCE_c_385_n N_VGND_c_1665_n 0.00469214f $X=0.87 $Y=0.2 $X2=0 $Y2=0
cc_363 N_SCE_c_384_n N_VGND_c_1667_n 0.0380833f $X=2.265 $Y=0.2 $X2=0 $Y2=0
cc_364 N_SCE_c_384_n N_VGND_c_1680_n 0.0552899f $X=2.265 $Y=0.2 $X2=0 $Y2=0
cc_365 N_SCE_c_385_n N_VGND_c_1680_n 0.00952178f $X=0.87 $Y=0.2 $X2=0 $Y2=0
cc_366 N_SCD_M1026_g N_CLK_M1028_g 0.0196032f $X=2.7 $Y=0.825 $X2=0 $Y2=0
cc_367 N_SCD_M1001_g N_CLK_c_497_n 0.0412554f $X=2.665 $Y=2.775 $X2=0 $Y2=0
cc_368 SCD N_CLK_c_497_n 3.65396e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_369 N_SCD_c_453_n N_CLK_c_497_n 0.0196032f $X=2.61 $Y=1.56 $X2=0 $Y2=0
cc_370 N_SCD_M1001_g N_A_641_123#_c_573_n 3.85276e-19 $X=2.665 $Y=2.775 $X2=0
+ $Y2=0
cc_371 N_SCD_M1001_g N_VPWR_c_1331_n 0.00617328f $X=2.665 $Y=2.775 $X2=0 $Y2=0
cc_372 N_SCD_M1001_g N_VPWR_c_1337_n 0.00502699f $X=2.665 $Y=2.775 $X2=0 $Y2=0
cc_373 N_SCD_M1001_g N_VPWR_c_1329_n 0.00630632f $X=2.665 $Y=2.775 $X2=0 $Y2=0
cc_374 N_SCD_M1001_g N_A_359_123#_c_1497_n 0.00940762f $X=2.665 $Y=2.775 $X2=0
+ $Y2=0
cc_375 N_SCD_M1026_g N_A_359_123#_c_1485_n 0.0156963f $X=2.7 $Y=0.825 $X2=0
+ $Y2=0
cc_376 SCD N_A_359_123#_c_1485_n 0.0440147f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_377 N_SCD_c_453_n N_A_359_123#_c_1485_n 0.0041462f $X=2.61 $Y=1.56 $X2=0
+ $Y2=0
cc_378 SCD N_A_359_123#_c_1486_n 0.0159602f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_379 N_SCD_M1001_g N_A_359_123#_c_1500_n 0.00402884f $X=2.665 $Y=2.775 $X2=0
+ $Y2=0
cc_380 N_SCD_M1001_g N_A_359_123#_c_1487_n 0.00598705f $X=2.665 $Y=2.775 $X2=0
+ $Y2=0
cc_381 N_SCD_M1026_g N_A_359_123#_c_1487_n 0.00615431f $X=2.7 $Y=0.825 $X2=0
+ $Y2=0
cc_382 SCD N_A_359_123#_c_1487_n 0.0304109f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_383 N_SCD_M1001_g N_A_359_123#_c_1502_n 0.00394335f $X=2.665 $Y=2.775 $X2=0
+ $Y2=0
cc_384 SCD N_A_359_123#_c_1502_n 0.00130215f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_385 N_SCD_M1001_g N_A_359_123#_c_1492_n 0.0165498f $X=2.665 $Y=2.775 $X2=0
+ $Y2=0
cc_386 SCD N_A_359_123#_c_1492_n 0.0101405f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_387 N_SCD_c_453_n N_A_359_123#_c_1492_n 0.0018791f $X=2.61 $Y=1.56 $X2=0
+ $Y2=0
cc_388 N_SCD_M1026_g N_VGND_c_1658_n 0.00930578f $X=2.7 $Y=0.825 $X2=0 $Y2=0
cc_389 N_SCD_M1026_g N_VGND_c_1667_n 0.00349617f $X=2.7 $Y=0.825 $X2=0 $Y2=0
cc_390 N_SCD_M1026_g N_VGND_c_1680_n 0.00396651f $X=2.7 $Y=0.825 $X2=0 $Y2=0
cc_391 CLK N_A_641_123#_c_540_n 0.00220196f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_392 N_CLK_c_497_n N_A_641_123#_c_540_n 0.00588667f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_393 CLK N_A_641_123#_c_544_n 9.50146e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_394 N_CLK_c_497_n N_A_641_123#_c_544_n 0.00645593f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_395 N_CLK_M1028_g N_A_641_123#_c_548_n 0.00630216f $X=3.13 $Y=0.825 $X2=0
+ $Y2=0
cc_396 CLK N_A_641_123#_c_548_n 0.0357742f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_397 N_CLK_c_497_n N_A_641_123#_c_548_n 0.00154949f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_398 CLK N_A_641_123#_c_564_n 0.0133383f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_399 N_CLK_M1028_g N_A_641_123#_c_550_n 0.00276464f $X=3.13 $Y=0.825 $X2=0
+ $Y2=0
cc_400 N_CLK_M1031_g N_A_641_123#_c_550_n 0.00443071f $X=3.13 $Y=2.775 $X2=0
+ $Y2=0
cc_401 CLK N_A_641_123#_c_550_n 0.0808058f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_402 N_CLK_c_497_n N_A_641_123#_c_550_n 0.00185323f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_403 N_CLK_M1031_g N_A_641_123#_c_573_n 0.010925f $X=3.13 $Y=2.775 $X2=0 $Y2=0
cc_404 CLK N_A_641_123#_c_573_n 0.0159896f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_405 N_CLK_c_497_n N_A_641_123#_c_573_n 0.00112268f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_406 N_CLK_M1028_g N_A_641_123#_c_554_n 0.0039874f $X=3.13 $Y=0.825 $X2=0
+ $Y2=0
cc_407 N_CLK_M1031_g N_VPWR_c_1331_n 0.00320608f $X=3.13 $Y=2.775 $X2=0 $Y2=0
cc_408 N_CLK_M1031_g N_VPWR_c_1332_n 0.00225841f $X=3.13 $Y=2.775 $X2=0 $Y2=0
cc_409 N_CLK_M1031_g N_VPWR_c_1339_n 0.0054895f $X=3.13 $Y=2.775 $X2=0 $Y2=0
cc_410 N_CLK_M1031_g N_VPWR_c_1329_n 0.0112887f $X=3.13 $Y=2.775 $X2=0 $Y2=0
cc_411 N_CLK_M1028_g N_A_359_123#_c_1485_n 0.00918705f $X=3.13 $Y=0.825 $X2=0
+ $Y2=0
cc_412 CLK N_A_359_123#_c_1485_n 0.00199151f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_413 N_CLK_M1031_g N_A_359_123#_c_1500_n 5.39157e-19 $X=3.13 $Y=2.775 $X2=0
+ $Y2=0
cc_414 N_CLK_M1031_g N_A_359_123#_c_1487_n 0.00614136f $X=3.13 $Y=2.775 $X2=0
+ $Y2=0
cc_415 CLK N_A_359_123#_c_1487_n 0.064155f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_416 N_CLK_c_497_n N_A_359_123#_c_1487_n 0.0155824f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_417 N_CLK_M1031_g N_A_359_123#_c_1491_n 0.014174f $X=3.13 $Y=2.775 $X2=0
+ $Y2=0
cc_418 CLK N_A_359_123#_c_1491_n 0.00520534f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_419 N_CLK_c_497_n N_A_359_123#_c_1491_n 0.00118538f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_420 N_CLK_M1031_g N_A_359_123#_c_1502_n 4.19988e-19 $X=3.13 $Y=2.775 $X2=0
+ $Y2=0
cc_421 N_CLK_M1031_g N_A_359_123#_c_1492_n 0.0111984f $X=3.13 $Y=2.775 $X2=0
+ $Y2=0
cc_422 N_CLK_M1028_g N_VGND_c_1658_n 0.0163945f $X=3.13 $Y=0.825 $X2=0 $Y2=0
cc_423 N_CLK_M1028_g N_VGND_c_1659_n 0.00311696f $X=3.13 $Y=0.825 $X2=0 $Y2=0
cc_424 N_CLK_M1028_g N_VGND_c_1671_n 0.00349617f $X=3.13 $Y=0.825 $X2=0 $Y2=0
cc_425 N_CLK_M1028_g N_VGND_c_1680_n 0.00396651f $X=3.13 $Y=0.825 $X2=0 $Y2=0
cc_426 N_A_641_123#_c_566_n N_A_850_51#_M1003_d 0.00282402f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_427 N_A_641_123#_c_540_n N_A_850_51#_c_798_n 0.00614054f $X=4.175 $Y=2.145
+ $X2=0 $Y2=0
cc_428 N_A_641_123#_c_550_n N_A_850_51#_c_798_n 6.15096e-19 $X=4.082 $Y=2.3
+ $X2=0 $Y2=0
cc_429 N_A_641_123#_M1022_g N_A_850_51#_c_799_n 0.0146391f $X=5.92 $Y=2.455
+ $X2=0 $Y2=0
cc_430 N_A_641_123#_c_546_n N_A_850_51#_c_799_n 0.0194792f $X=5.265 $Y=1.68
+ $X2=0 $Y2=0
cc_431 N_A_641_123#_c_566_n N_A_850_51#_c_799_n 0.00147063f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_432 N_A_641_123#_c_568_n N_A_850_51#_c_799_n 2.81149e-19 $X=5.96 $Y=2.635
+ $X2=0 $Y2=0
cc_433 N_A_641_123#_c_561_n N_A_850_51#_c_800_n 0.00304182f $X=4.35 $Y=2.22
+ $X2=0 $Y2=0
cc_434 N_A_641_123#_c_566_n N_A_850_51#_c_800_n 0.0039407f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_435 N_A_641_123#_c_566_n N_A_850_51#_c_801_n 0.0070131f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_436 N_A_641_123#_c_576_n N_A_850_51#_c_801_n 0.00234301f $X=5.96 $Y=2.72
+ $X2=0 $Y2=0
cc_437 N_A_641_123#_M1009_g N_A_850_51#_c_780_n 0.0104325f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_438 N_A_641_123#_c_547_n N_A_850_51#_c_780_n 0.00501378f $X=5.845 $Y=1.68
+ $X2=0 $Y2=0
cc_439 N_A_641_123#_c_552_n N_A_850_51#_c_781_n 0.00424292f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_440 N_A_641_123#_c_553_n N_A_850_51#_c_781_n 9.69285e-19 $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_441 N_A_641_123#_c_556_n N_A_850_51#_c_781_n 0.00379412f $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_442 N_A_641_123#_c_551_n N_A_850_51#_c_782_n 0.003696f $X=7.89 $Y=1.825 $X2=0
+ $Y2=0
cc_443 N_A_641_123#_c_553_n N_A_850_51#_c_782_n 0.00456034f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_444 N_A_641_123#_c_556_n N_A_850_51#_c_782_n 0.0185756f $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_445 N_A_641_123#_c_571_n N_A_850_51#_c_783_n 0.00309098f $X=7.805 $Y=1.915
+ $X2=0 $Y2=0
cc_446 N_A_641_123#_c_551_n N_A_850_51#_c_783_n 0.00134611f $X=7.89 $Y=1.825
+ $X2=0 $Y2=0
cc_447 N_A_641_123#_c_556_n N_A_850_51#_c_783_n 0.00199816f $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_448 N_A_641_123#_M1023_g N_A_850_51#_M1032_g 0.0110277f $X=7.3 $Y=2.665 $X2=0
+ $Y2=0
cc_449 N_A_641_123#_c_570_n N_A_850_51#_M1032_g 0.00424342f $X=7.515 $Y=2.635
+ $X2=0 $Y2=0
cc_450 N_A_641_123#_c_571_n N_A_850_51#_M1032_g 0.00186371f $X=7.805 $Y=1.915
+ $X2=0 $Y2=0
cc_451 N_A_641_123#_c_551_n N_A_850_51#_M1032_g 0.00611811f $X=7.89 $Y=1.825
+ $X2=0 $Y2=0
cc_452 N_A_641_123#_c_577_n N_A_850_51#_M1032_g 0.00797994f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_453 N_A_641_123#_c_545_n N_A_850_51#_c_803_n 0.0183341f $X=4.085 $Y=1.455
+ $X2=0 $Y2=0
cc_454 N_A_641_123#_c_546_n N_A_850_51#_c_803_n 0.0120861f $X=5.265 $Y=1.68
+ $X2=0 $Y2=0
cc_455 N_A_641_123#_M1009_g N_A_850_51#_c_785_n 2.54929e-19 $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_456 N_A_641_123#_c_544_n N_A_850_51#_c_785_n 0.00185667f $X=4.085 $Y=1.29
+ $X2=0 $Y2=0
cc_457 N_A_641_123#_c_545_n N_A_850_51#_c_786_n 0.00185667f $X=4.085 $Y=1.455
+ $X2=0 $Y2=0
cc_458 N_A_641_123#_c_561_n N_A_850_51#_c_786_n 0.00515468f $X=4.35 $Y=2.22
+ $X2=0 $Y2=0
cc_459 N_A_641_123#_c_546_n N_A_850_51#_c_786_n 2.54929e-19 $X=5.265 $Y=1.68
+ $X2=0 $Y2=0
cc_460 N_A_641_123#_c_630_p N_A_850_51#_c_786_n 0.00861606f $X=4.215 $Y=2.895
+ $X2=0 $Y2=0
cc_461 N_A_641_123#_c_566_n N_A_850_51#_c_786_n 0.0196291f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_462 N_A_641_123#_c_574_n N_A_850_51#_c_786_n 0.0109651f $X=4.082 $Y=2.385
+ $X2=0 $Y2=0
cc_463 N_A_641_123#_M1009_g N_A_850_51#_c_787_n 0.0120861f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_464 N_A_641_123#_c_544_n N_A_850_51#_c_787_n 0.0183341f $X=4.085 $Y=1.29
+ $X2=0 $Y2=0
cc_465 N_A_641_123#_c_550_n N_A_850_51#_c_787_n 0.00227118f $X=4.082 $Y=2.3
+ $X2=0 $Y2=0
cc_466 N_A_641_123#_M1009_g N_A_850_51#_c_788_n 0.0071049f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_467 N_A_641_123#_M1009_g N_A_850_51#_c_789_n 0.00133275f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_468 N_A_641_123#_M1034_g N_A_850_51#_c_791_n 0.00193902f $X=8.275 $Y=0.515
+ $X2=0 $Y2=0
cc_469 N_A_641_123#_M1034_g N_A_850_51#_c_792_n 0.00278883f $X=8.275 $Y=0.515
+ $X2=0 $Y2=0
cc_470 N_A_641_123#_c_571_n N_A_850_51#_c_792_n 0.00501903f $X=7.805 $Y=1.915
+ $X2=0 $Y2=0
cc_471 N_A_641_123#_c_552_n N_A_850_51#_c_792_n 0.0226766f $X=8.25 $Y=1.02 $X2=0
+ $Y2=0
cc_472 N_A_641_123#_c_553_n N_A_850_51#_c_792_n 2.79484e-19 $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_473 N_A_641_123#_M1034_g N_A_850_51#_c_793_n 7.32804e-19 $X=8.275 $Y=0.515
+ $X2=0 $Y2=0
cc_474 N_A_641_123#_c_571_n N_A_850_51#_c_793_n 7.76658e-19 $X=7.805 $Y=1.915
+ $X2=0 $Y2=0
cc_475 N_A_641_123#_c_552_n N_A_850_51#_c_793_n 0.00208842f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_476 N_A_641_123#_c_553_n N_A_850_51#_c_793_n 0.0192486f $X=8.25 $Y=1.02 $X2=0
+ $Y2=0
cc_477 N_A_641_123#_c_577_n N_A_850_51#_c_793_n 0.00160745f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_478 N_A_641_123#_c_578_n N_A_850_51#_c_793_n 3.70564e-19 $X=7.6 $Y=1.93 $X2=0
+ $Y2=0
cc_479 N_A_641_123#_c_556_n N_A_850_51#_c_793_n 8.02523e-19 $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_480 N_A_641_123#_M1009_g N_A_850_51#_c_794_n 0.00277854f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_481 N_A_641_123#_M1009_g N_A_850_51#_c_795_n 0.00288031f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_482 N_A_641_123#_c_543_n N_A_850_51#_c_795_n 0.00550678f $X=4.085 $Y=0.785
+ $X2=0 $Y2=0
cc_483 N_A_641_123#_c_549_n N_A_850_51#_c_795_n 0.0200327f $X=4.082 $Y=1.02
+ $X2=0 $Y2=0
cc_484 N_A_641_123#_c_550_n N_A_850_51#_c_795_n 0.106175f $X=4.082 $Y=2.3 $X2=0
+ $Y2=0
cc_485 N_A_641_123#_c_554_n N_A_850_51#_c_795_n 0.00185667f $X=4.085 $Y=0.95
+ $X2=0 $Y2=0
cc_486 N_A_641_123#_M1034_g N_A_850_51#_c_797_n 0.00885502f $X=8.275 $Y=0.515
+ $X2=0 $Y2=0
cc_487 N_A_641_123#_c_569_n N_A_1203_99#_M1002_d 0.00427471f $X=7.43 $Y=2.72
+ $X2=0 $Y2=0
cc_488 N_A_641_123#_c_547_n N_A_1203_99#_c_956_n 0.0391269f $X=5.845 $Y=1.68
+ $X2=0 $Y2=0
cc_489 N_A_641_123#_c_555_n N_A_1203_99#_c_956_n 0.00272182f $X=5.96 $Y=1.68
+ $X2=0 $Y2=0
cc_490 N_A_641_123#_c_568_n N_A_1203_99#_c_957_n 0.00571572f $X=5.96 $Y=2.635
+ $X2=0 $Y2=0
cc_491 N_A_641_123#_c_569_n N_A_1203_99#_M1021_g 0.0121725f $X=7.43 $Y=2.72
+ $X2=0 $Y2=0
cc_492 N_A_641_123#_M1022_g N_A_1203_99#_c_964_n 0.0391269f $X=5.92 $Y=2.455
+ $X2=0 $Y2=0
cc_493 N_A_641_123#_c_569_n N_A_1203_99#_c_964_n 0.00361875f $X=7.43 $Y=2.72
+ $X2=0 $Y2=0
cc_494 N_A_641_123#_M1022_g N_A_1203_99#_c_958_n 2.50877e-19 $X=5.92 $Y=2.455
+ $X2=0 $Y2=0
cc_495 N_A_641_123#_M1023_g N_A_1203_99#_c_958_n 0.00421789f $X=7.3 $Y=2.665
+ $X2=0 $Y2=0
cc_496 N_A_641_123#_c_547_n N_A_1203_99#_c_958_n 3.51999e-19 $X=5.845 $Y=1.68
+ $X2=0 $Y2=0
cc_497 N_A_641_123#_c_568_n N_A_1203_99#_c_958_n 0.0174812f $X=5.96 $Y=2.635
+ $X2=0 $Y2=0
cc_498 N_A_641_123#_c_569_n N_A_1203_99#_c_958_n 0.0361354f $X=7.43 $Y=2.72
+ $X2=0 $Y2=0
cc_499 N_A_641_123#_c_570_n N_A_1203_99#_c_958_n 0.0164028f $X=7.515 $Y=2.635
+ $X2=0 $Y2=0
cc_500 N_A_641_123#_c_555_n N_A_1203_99#_c_958_n 0.0264688f $X=5.96 $Y=1.68
+ $X2=0 $Y2=0
cc_501 N_A_641_123#_c_577_n N_A_1203_99#_c_958_n 0.00482302f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_502 N_A_641_123#_c_578_n N_A_1203_99#_c_958_n 0.017672f $X=7.6 $Y=1.93 $X2=0
+ $Y2=0
cc_503 N_A_641_123#_c_577_n N_A_1203_99#_c_959_n 0.00660669f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_504 N_A_641_123#_c_578_n N_A_1203_99#_c_959_n 0.0142329f $X=7.6 $Y=1.93 $X2=0
+ $Y2=0
cc_505 N_A_641_123#_c_556_n N_A_1203_99#_c_959_n 0.00887887f $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_506 N_A_641_123#_c_552_n N_A_1203_99#_c_960_n 0.00646421f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_507 N_A_641_123#_c_556_n N_A_1203_99#_c_960_n 0.00573523f $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_508 N_A_641_123#_c_569_n N_A_1053_125#_M1002_g 0.0136578f $X=7.43 $Y=2.72
+ $X2=0 $Y2=0
cc_509 N_A_641_123#_c_577_n N_A_1053_125#_M1002_g 0.0523762f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_510 N_A_641_123#_c_547_n N_A_1053_125#_c_1023_n 0.0105744f $X=5.845 $Y=1.68
+ $X2=0 $Y2=0
cc_511 N_A_641_123#_c_555_n N_A_1053_125#_c_1023_n 0.0221995f $X=5.96 $Y=1.68
+ $X2=0 $Y2=0
cc_512 N_A_641_123#_M1009_g N_A_1053_125#_c_1024_n 0.00395198f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_513 N_A_641_123#_c_547_n N_A_1053_125#_c_1024_n 0.0017469f $X=5.845 $Y=1.68
+ $X2=0 $Y2=0
cc_514 N_A_641_123#_M1022_g N_A_1053_125#_c_1028_n 0.00413503f $X=5.92 $Y=2.455
+ $X2=0 $Y2=0
cc_515 N_A_641_123#_c_547_n N_A_1053_125#_c_1028_n 0.00557939f $X=5.845 $Y=1.68
+ $X2=0 $Y2=0
cc_516 N_A_641_123#_c_566_n N_A_1053_125#_c_1028_n 0.0240254f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_517 N_A_641_123#_c_568_n N_A_1053_125#_c_1028_n 0.0371267f $X=5.96 $Y=2.635
+ $X2=0 $Y2=0
cc_518 N_A_641_123#_M1009_g N_A_1053_125#_c_1025_n 0.00448753f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_519 N_A_641_123#_M1022_g N_A_1053_125#_c_1025_n 0.00495365f $X=5.92 $Y=2.455
+ $X2=0 $Y2=0
cc_520 N_A_641_123#_c_547_n N_A_1053_125#_c_1025_n 0.0232817f $X=5.845 $Y=1.68
+ $X2=0 $Y2=0
cc_521 N_A_641_123#_c_568_n N_A_1053_125#_c_1025_n 0.0164515f $X=5.96 $Y=2.635
+ $X2=0 $Y2=0
cc_522 N_A_641_123#_c_555_n N_A_1053_125#_c_1025_n 0.023673f $X=5.96 $Y=1.68
+ $X2=0 $Y2=0
cc_523 N_A_641_123#_M1034_g N_A_1673_409#_M1029_g 0.0309909f $X=8.275 $Y=0.515
+ $X2=0 $Y2=0
cc_524 N_A_641_123#_c_552_n N_A_1673_409#_M1029_g 0.00191106f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_525 N_A_641_123#_c_553_n N_A_1673_409#_M1029_g 0.0203555f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_526 N_A_641_123#_c_569_n N_A_1475_449#_M1023_d 0.00468341f $X=7.43 $Y=2.72
+ $X2=0 $Y2=0
cc_527 N_A_641_123#_c_570_n N_A_1475_449#_M1023_d 0.00781468f $X=7.515 $Y=2.635
+ $X2=0 $Y2=0
cc_528 N_A_641_123#_M1023_g N_A_1475_449#_c_1247_n 0.00291744f $X=7.3 $Y=2.665
+ $X2=0 $Y2=0
cc_529 N_A_641_123#_c_569_n N_A_1475_449#_c_1247_n 0.0151f $X=7.43 $Y=2.72 $X2=0
+ $Y2=0
cc_530 N_A_641_123#_c_570_n N_A_1475_449#_c_1247_n 0.00428495f $X=7.515 $Y=2.635
+ $X2=0 $Y2=0
cc_531 N_A_641_123#_c_571_n N_A_1475_449#_c_1247_n 0.00677369f $X=7.805 $Y=1.915
+ $X2=0 $Y2=0
cc_532 N_A_641_123#_M1034_g N_A_1475_449#_c_1251_n 0.0126794f $X=8.275 $Y=0.515
+ $X2=0 $Y2=0
cc_533 N_A_641_123#_c_552_n N_A_1475_449#_c_1251_n 0.0252517f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_534 N_A_641_123#_c_553_n N_A_1475_449#_c_1251_n 0.00215414f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_535 N_A_641_123#_c_556_n N_A_1475_449#_c_1251_n 3.20559e-19 $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_536 N_A_641_123#_c_570_n N_A_1475_449#_c_1240_n 0.0164782f $X=7.515 $Y=2.635
+ $X2=0 $Y2=0
cc_537 N_A_641_123#_c_571_n N_A_1475_449#_c_1240_n 0.0113432f $X=7.805 $Y=1.915
+ $X2=0 $Y2=0
cc_538 N_A_641_123#_c_578_n N_A_1475_449#_c_1240_n 8.87036e-19 $X=7.6 $Y=1.93
+ $X2=0 $Y2=0
cc_539 N_A_641_123#_c_553_n N_A_1475_449#_c_1241_n 0.00220488f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_540 N_A_641_123#_c_556_n N_A_1475_449#_c_1241_n 6.91831e-19 $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_541 N_A_641_123#_c_571_n N_A_1475_449#_c_1242_n 0.00336326f $X=7.805 $Y=1.915
+ $X2=0 $Y2=0
cc_542 N_A_641_123#_c_551_n N_A_1475_449#_c_1242_n 0.00971438f $X=7.89 $Y=1.825
+ $X2=0 $Y2=0
cc_543 N_A_641_123#_c_553_n N_A_1475_449#_c_1242_n 6.6652e-19 $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_544 N_A_641_123#_c_556_n N_A_1475_449#_c_1242_n 0.0152576f $X=8.07 $Y=1.515
+ $X2=0 $Y2=0
cc_545 N_A_641_123#_M1034_g N_A_1475_449#_c_1233_n 0.00371465f $X=8.275 $Y=0.515
+ $X2=0 $Y2=0
cc_546 N_A_641_123#_c_552_n N_A_1475_449#_c_1233_n 0.0238758f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_547 N_A_641_123#_c_553_n N_A_1475_449#_c_1233_n 0.00204684f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_548 N_A_641_123#_c_551_n N_A_1475_449#_c_1234_n 0.0058817f $X=7.89 $Y=1.825
+ $X2=0 $Y2=0
cc_549 N_A_641_123#_c_552_n N_A_1475_449#_c_1237_n 0.0287072f $X=8.25 $Y=1.02
+ $X2=0 $Y2=0
cc_550 N_A_641_123#_c_564_n N_VPWR_M1003_s 0.00102363f $X=3.865 $Y=2.385 $X2=0
+ $Y2=0
cc_551 N_A_641_123#_c_630_p N_VPWR_M1003_s 0.00585449f $X=4.215 $Y=2.895 $X2=0
+ $Y2=0
cc_552 N_A_641_123#_c_567_n N_VPWR_M1003_s 0.00166402f $X=4.3 $Y=2.98 $X2=0
+ $Y2=0
cc_553 N_A_641_123#_c_574_n N_VPWR_M1003_s 0.00356706f $X=4.082 $Y=2.385 $X2=0
+ $Y2=0
cc_554 N_A_641_123#_c_569_n N_VPWR_M1021_d 0.00966977f $X=7.43 $Y=2.72 $X2=0
+ $Y2=0
cc_555 N_A_641_123#_c_558_n N_VPWR_c_1332_n 0.00476612f $X=4.35 $Y=2.295 $X2=0
+ $Y2=0
cc_556 N_A_641_123#_c_564_n N_VPWR_c_1332_n 0.0117026f $X=3.865 $Y=2.385 $X2=0
+ $Y2=0
cc_557 N_A_641_123#_c_630_p N_VPWR_c_1332_n 0.0190935f $X=4.215 $Y=2.895 $X2=0
+ $Y2=0
cc_558 N_A_641_123#_c_567_n N_VPWR_c_1332_n 0.0143027f $X=4.3 $Y=2.98 $X2=0
+ $Y2=0
cc_559 N_A_641_123#_c_573_n N_VPWR_c_1332_n 0.0328737f $X=3.345 $Y=2.61 $X2=0
+ $Y2=0
cc_560 N_A_641_123#_c_574_n N_VPWR_c_1332_n 0.00680349f $X=4.082 $Y=2.385 $X2=0
+ $Y2=0
cc_561 N_A_641_123#_c_573_n N_VPWR_c_1339_n 0.0209566f $X=3.345 $Y=2.61 $X2=0
+ $Y2=0
cc_562 N_A_641_123#_c_558_n N_VPWR_c_1344_n 0.00327695f $X=4.35 $Y=2.295 $X2=0
+ $Y2=0
cc_563 N_A_641_123#_M1022_g N_VPWR_c_1344_n 4.48664e-19 $X=5.92 $Y=2.455 $X2=0
+ $Y2=0
cc_564 N_A_641_123#_c_566_n N_VPWR_c_1344_n 0.095117f $X=5.875 $Y=2.98 $X2=0
+ $Y2=0
cc_565 N_A_641_123#_c_567_n N_VPWR_c_1344_n 0.0113451f $X=4.3 $Y=2.98 $X2=0
+ $Y2=0
cc_566 N_A_641_123#_c_569_n N_VPWR_c_1344_n 0.00857039f $X=7.43 $Y=2.72 $X2=0
+ $Y2=0
cc_567 N_A_641_123#_c_576_n N_VPWR_c_1344_n 0.0113273f $X=5.96 $Y=2.72 $X2=0
+ $Y2=0
cc_568 N_A_641_123#_M1023_g N_VPWR_c_1345_n 0.00400062f $X=7.3 $Y=2.665 $X2=0
+ $Y2=0
cc_569 N_A_641_123#_c_569_n N_VPWR_c_1345_n 0.0173604f $X=7.43 $Y=2.72 $X2=0
+ $Y2=0
cc_570 N_A_641_123#_c_569_n N_VPWR_c_1349_n 0.0240258f $X=7.43 $Y=2.72 $X2=0
+ $Y2=0
cc_571 N_A_641_123#_c_576_n N_VPWR_c_1349_n 0.00420802f $X=5.96 $Y=2.72 $X2=0
+ $Y2=0
cc_572 N_A_641_123#_M1031_d N_VPWR_c_1329_n 0.00215158f $X=3.205 $Y=2.455 $X2=0
+ $Y2=0
cc_573 N_A_641_123#_c_558_n N_VPWR_c_1329_n 0.00667022f $X=4.35 $Y=2.295 $X2=0
+ $Y2=0
cc_574 N_A_641_123#_M1023_g N_VPWR_c_1329_n 0.00698731f $X=7.3 $Y=2.665 $X2=0
+ $Y2=0
cc_575 N_A_641_123#_c_564_n N_VPWR_c_1329_n 0.00425342f $X=3.865 $Y=2.385 $X2=0
+ $Y2=0
cc_576 N_A_641_123#_c_566_n N_VPWR_c_1329_n 0.0582868f $X=5.875 $Y=2.98 $X2=0
+ $Y2=0
cc_577 N_A_641_123#_c_567_n N_VPWR_c_1329_n 0.00645785f $X=4.3 $Y=2.98 $X2=0
+ $Y2=0
cc_578 N_A_641_123#_c_569_n N_VPWR_c_1329_n 0.0387536f $X=7.43 $Y=2.72 $X2=0
+ $Y2=0
cc_579 N_A_641_123#_c_573_n N_VPWR_c_1329_n 0.0125409f $X=3.345 $Y=2.61 $X2=0
+ $Y2=0
cc_580 N_A_641_123#_c_574_n N_VPWR_c_1329_n 0.00367988f $X=4.082 $Y=2.385 $X2=0
+ $Y2=0
cc_581 N_A_641_123#_c_576_n N_VPWR_c_1329_n 0.00650045f $X=5.96 $Y=2.72 $X2=0
+ $Y2=0
cc_582 N_A_641_123#_c_573_n N_A_359_123#_c_1497_n 6.285e-19 $X=3.345 $Y=2.61
+ $X2=0 $Y2=0
cc_583 N_A_641_123#_c_573_n N_A_359_123#_c_1500_n 0.00359097f $X=3.345 $Y=2.61
+ $X2=0 $Y2=0
cc_584 N_A_641_123#_M1009_g N_A_359_123#_c_1488_n 0.00388235f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_585 N_A_641_123#_M1031_d N_A_359_123#_c_1491_n 9.59932e-19 $X=3.205 $Y=2.455
+ $X2=0 $Y2=0
cc_586 N_A_641_123#_c_558_n N_A_359_123#_c_1491_n 0.00713861f $X=4.35 $Y=2.295
+ $X2=0 $Y2=0
cc_587 N_A_641_123#_c_564_n N_A_359_123#_c_1491_n 0.0181133f $X=3.865 $Y=2.385
+ $X2=0 $Y2=0
cc_588 N_A_641_123#_c_630_p N_A_359_123#_c_1491_n 0.00905213f $X=4.215 $Y=2.895
+ $X2=0 $Y2=0
cc_589 N_A_641_123#_c_566_n N_A_359_123#_c_1491_n 0.0115627f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_590 N_A_641_123#_c_573_n N_A_359_123#_c_1491_n 0.0234074f $X=3.345 $Y=2.61
+ $X2=0 $Y2=0
cc_591 N_A_641_123#_c_574_n N_A_359_123#_c_1491_n 0.0287112f $X=4.082 $Y=2.385
+ $X2=0 $Y2=0
cc_592 N_A_641_123#_c_573_n N_A_359_123#_c_1502_n 0.00112147f $X=3.345 $Y=2.61
+ $X2=0 $Y2=0
cc_593 N_A_641_123#_c_573_n N_A_359_123#_c_1492_n 0.00740679f $X=3.345 $Y=2.61
+ $X2=0 $Y2=0
cc_594 N_A_641_123#_c_566_n N_A_359_123#_c_1493_n 0.00255095f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_595 N_A_641_123#_c_566_n N_A_359_123#_c_1494_n 0.0118419f $X=5.875 $Y=2.98
+ $X2=0 $Y2=0
cc_596 N_A_641_123#_M1009_g N_A_359_123#_c_1489_n 0.0125014f $X=5.19 $Y=0.835
+ $X2=0 $Y2=0
cc_597 N_A_641_123#_c_546_n N_A_359_123#_c_1489_n 0.00934946f $X=5.265 $Y=1.68
+ $X2=0 $Y2=0
cc_598 N_A_641_123#_c_569_n A_1199_449# 0.00366293f $X=7.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.245
cc_599 N_A_641_123#_c_548_n N_VGND_c_1658_n 0.00660981f $X=3.865 $Y=0.902 $X2=0
+ $Y2=0
cc_600 N_A_641_123#_c_543_n N_VGND_c_1659_n 0.0103434f $X=4.085 $Y=0.785 $X2=0
+ $Y2=0
cc_601 N_A_641_123#_c_548_n N_VGND_c_1659_n 0.00571776f $X=3.865 $Y=0.902 $X2=0
+ $Y2=0
cc_602 N_A_641_123#_c_549_n N_VGND_c_1659_n 0.0195819f $X=4.082 $Y=1.02 $X2=0
+ $Y2=0
cc_603 N_A_641_123#_c_554_n N_VGND_c_1659_n 0.00123408f $X=4.085 $Y=0.95 $X2=0
+ $Y2=0
cc_604 N_A_641_123#_c_543_n N_VGND_c_1672_n 0.00469214f $X=4.085 $Y=0.785 $X2=0
+ $Y2=0
cc_605 N_A_641_123#_M1034_g N_VGND_c_1673_n 0.00329012f $X=8.275 $Y=0.515 $X2=0
+ $Y2=0
cc_606 N_A_641_123#_M1034_g N_VGND_c_1680_n 0.00496803f $X=8.275 $Y=0.515 $X2=0
+ $Y2=0
cc_607 N_A_641_123#_c_543_n N_VGND_c_1680_n 0.00559969f $X=4.085 $Y=0.785 $X2=0
+ $Y2=0
cc_608 N_A_641_123#_c_548_n N_VGND_c_1680_n 0.0197022f $X=3.865 $Y=0.902 $X2=0
+ $Y2=0
cc_609 N_A_641_123#_c_549_n N_VGND_c_1680_n 0.0070574f $X=4.082 $Y=1.02 $X2=0
+ $Y2=0
cc_610 N_A_850_51#_c_791_n N_A_1203_99#_M1019_d 0.00415348f $X=7.615 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_611 N_A_850_51#_c_780_n N_A_1203_99#_c_955_n 0.0265128f $X=5.64 $Y=0.515
+ $X2=0 $Y2=0
cc_612 N_A_850_51#_c_788_n N_A_1203_99#_c_955_n 0.00154532f $X=5.72 $Y=0.375
+ $X2=0 $Y2=0
cc_613 N_A_850_51#_c_789_n N_A_1203_99#_c_955_n 0.00117589f $X=5.64 $Y=0.35
+ $X2=0 $Y2=0
cc_614 N_A_850_51#_c_790_n N_A_1203_99#_c_955_n 0.012473f $X=6.765 $Y=0.64 $X2=0
+ $Y2=0
cc_615 N_A_850_51#_c_796_n N_A_1203_99#_c_955_n 0.00166789f $X=6.85 $Y=0.34
+ $X2=0 $Y2=0
cc_616 N_A_850_51#_c_790_n N_A_1203_99#_c_956_n 8.15688e-19 $X=6.765 $Y=0.64
+ $X2=0 $Y2=0
cc_617 N_A_850_51#_c_783_n N_A_1203_99#_c_959_n 0.00176324f $X=7.845 $Y=1.47
+ $X2=0 $Y2=0
cc_618 N_A_850_51#_c_781_n N_A_1203_99#_c_960_n 0.00426973f $X=7.77 $Y=1.395
+ $X2=0 $Y2=0
cc_619 N_A_850_51#_c_793_n N_A_1203_99#_c_960_n 0.00247517f $X=7.71 $Y=1 $X2=0
+ $Y2=0
cc_620 N_A_850_51#_c_791_n N_A_1203_99#_c_961_n 0.0200016f $X=7.615 $Y=0.34
+ $X2=0 $Y2=0
cc_621 N_A_850_51#_c_792_n N_A_1203_99#_c_961_n 0.0418224f $X=7.71 $Y=1 $X2=0
+ $Y2=0
cc_622 N_A_850_51#_c_797_n N_A_1203_99#_c_961_n 0.00247517f $X=7.705 $Y=0.835
+ $X2=0 $Y2=0
cc_623 N_A_850_51#_c_791_n N_A_1053_125#_c_1022_n 0.0126943f $X=7.615 $Y=0.34
+ $X2=0 $Y2=0
cc_624 N_A_850_51#_c_792_n N_A_1053_125#_c_1022_n 6.69848e-19 $X=7.71 $Y=1 $X2=0
+ $Y2=0
cc_625 N_A_850_51#_c_796_n N_A_1053_125#_c_1022_n 0.00150242f $X=6.85 $Y=0.34
+ $X2=0 $Y2=0
cc_626 N_A_850_51#_c_797_n N_A_1053_125#_c_1022_n 0.0102804f $X=7.705 $Y=0.835
+ $X2=0 $Y2=0
cc_627 N_A_850_51#_c_780_n N_A_1053_125#_c_1049_n 3.22004e-19 $X=5.64 $Y=0.515
+ $X2=0 $Y2=0
cc_628 N_A_850_51#_c_788_n N_A_1053_125#_c_1049_n 0.0162761f $X=5.72 $Y=0.375
+ $X2=0 $Y2=0
cc_629 N_A_850_51#_c_789_n N_A_1053_125#_c_1049_n 0.00163585f $X=5.64 $Y=0.35
+ $X2=0 $Y2=0
cc_630 N_A_850_51#_c_780_n N_A_1053_125#_c_1023_n 0.00953803f $X=5.64 $Y=0.515
+ $X2=0 $Y2=0
cc_631 N_A_850_51#_c_788_n N_A_1053_125#_c_1023_n 0.0119281f $X=5.72 $Y=0.375
+ $X2=0 $Y2=0
cc_632 N_A_850_51#_c_789_n N_A_1053_125#_c_1023_n 7.36273e-19 $X=5.64 $Y=0.35
+ $X2=0 $Y2=0
cc_633 N_A_850_51#_c_790_n N_A_1053_125#_c_1023_n 0.0380759f $X=6.765 $Y=0.64
+ $X2=0 $Y2=0
cc_634 N_A_850_51#_c_791_n N_A_1053_125#_c_1023_n 0.00313622f $X=7.615 $Y=0.34
+ $X2=0 $Y2=0
cc_635 N_A_850_51#_c_796_n N_A_1053_125#_c_1023_n 0.00790791f $X=6.85 $Y=0.34
+ $X2=0 $Y2=0
cc_636 N_A_850_51#_c_801_n N_A_1053_125#_c_1028_n 0.0134575f $X=5.3 $Y=2.205
+ $X2=0 $Y2=0
cc_637 N_A_850_51#_c_786_n N_A_1053_125#_c_1028_n 0.00297682f $X=4.655 $Y=1.4
+ $X2=0 $Y2=0
cc_638 N_A_850_51#_c_799_n N_A_1053_125#_c_1025_n 0.0043405f $X=5.225 $Y=2.13
+ $X2=0 $Y2=0
cc_639 N_A_850_51#_c_801_n N_A_1053_125#_c_1025_n 4.05511e-19 $X=5.3 $Y=2.205
+ $X2=0 $Y2=0
cc_640 N_A_850_51#_c_781_n N_A_1053_125#_c_1026_n 0.00302817f $X=7.77 $Y=1.395
+ $X2=0 $Y2=0
cc_641 N_A_850_51#_c_793_n N_A_1053_125#_c_1026_n 0.0102804f $X=7.71 $Y=1 $X2=0
+ $Y2=0
cc_642 N_A_850_51#_c_796_n N_A_1053_125#_c_1026_n 0.0039543f $X=6.85 $Y=0.34
+ $X2=0 $Y2=0
cc_643 N_A_850_51#_c_782_n N_A_1673_409#_M1029_g 0.0129134f $X=8.005 $Y=1.47
+ $X2=0 $Y2=0
cc_644 N_A_850_51#_M1032_g N_A_1673_409#_c_1120_n 0.0590452f $X=8.08 $Y=2.745
+ $X2=0 $Y2=0
cc_645 N_A_850_51#_c_791_n N_A_1475_449#_M1033_d 0.0014369f $X=7.615 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_646 N_A_850_51#_c_792_n N_A_1475_449#_M1033_d 0.00299823f $X=7.71 $Y=1
+ $X2=-0.19 $Y2=-0.245
cc_647 N_A_850_51#_M1032_g N_A_1475_449#_c_1247_n 0.0155825f $X=8.08 $Y=2.745
+ $X2=0 $Y2=0
cc_648 N_A_850_51#_c_791_n N_A_1475_449#_c_1251_n 0.00715304f $X=7.615 $Y=0.34
+ $X2=0 $Y2=0
cc_649 N_A_850_51#_c_792_n N_A_1475_449#_c_1251_n 0.0203947f $X=7.71 $Y=1 $X2=0
+ $Y2=0
cc_650 N_A_850_51#_c_797_n N_A_1475_449#_c_1251_n 0.00117546f $X=7.705 $Y=0.835
+ $X2=0 $Y2=0
cc_651 N_A_850_51#_M1032_g N_A_1475_449#_c_1240_n 0.008252f $X=8.08 $Y=2.745
+ $X2=0 $Y2=0
cc_652 N_A_850_51#_M1032_g N_A_1475_449#_c_1242_n 0.00196662f $X=8.08 $Y=2.745
+ $X2=0 $Y2=0
cc_653 N_A_850_51#_c_782_n N_A_1475_449#_c_1234_n 0.00145598f $X=8.005 $Y=1.47
+ $X2=0 $Y2=0
cc_654 N_A_850_51#_c_782_n N_A_1475_449#_c_1237_n 3.63632e-19 $X=8.005 $Y=1.47
+ $X2=0 $Y2=0
cc_655 N_A_850_51#_M1032_g N_VPWR_c_1345_n 0.00298026f $X=8.08 $Y=2.745 $X2=0
+ $Y2=0
cc_656 N_A_850_51#_M1032_g N_VPWR_c_1350_n 0.00110585f $X=8.08 $Y=2.745 $X2=0
+ $Y2=0
cc_657 N_A_850_51#_M1032_g N_VPWR_c_1329_n 0.00544287f $X=8.08 $Y=2.745 $X2=0
+ $Y2=0
cc_658 N_A_850_51#_c_788_n N_A_359_123#_c_1488_n 0.0224409f $X=5.72 $Y=0.375
+ $X2=0 $Y2=0
cc_659 N_A_850_51#_c_795_n N_A_359_123#_c_1488_n 0.0263293f $X=4.61 $Y=1.235
+ $X2=0 $Y2=0
cc_660 N_A_850_51#_M1003_d N_A_359_123#_c_1491_n 4.60701e-19 $X=4.425 $Y=2.405
+ $X2=0 $Y2=0
cc_661 N_A_850_51#_c_800_n N_A_359_123#_c_1491_n 0.00363037f $X=4.82 $Y=2.13
+ $X2=0 $Y2=0
cc_662 N_A_850_51#_c_786_n N_A_359_123#_c_1491_n 0.0196122f $X=4.655 $Y=1.4
+ $X2=0 $Y2=0
cc_663 N_A_850_51#_c_799_n N_A_359_123#_c_1493_n 0.00149443f $X=5.225 $Y=2.13
+ $X2=0 $Y2=0
cc_664 N_A_850_51#_c_786_n N_A_359_123#_c_1493_n 0.00267659f $X=4.655 $Y=1.4
+ $X2=0 $Y2=0
cc_665 N_A_850_51#_c_799_n N_A_359_123#_c_1494_n 0.00140652f $X=5.225 $Y=2.13
+ $X2=0 $Y2=0
cc_666 N_A_850_51#_c_801_n N_A_359_123#_c_1494_n 4.52926e-19 $X=5.3 $Y=2.205
+ $X2=0 $Y2=0
cc_667 N_A_850_51#_c_786_n N_A_359_123#_c_1494_n 0.0522124f $X=4.655 $Y=1.4
+ $X2=0 $Y2=0
cc_668 N_A_850_51#_c_799_n N_A_359_123#_c_1489_n 0.0174266f $X=5.225 $Y=2.13
+ $X2=0 $Y2=0
cc_669 N_A_850_51#_c_801_n N_A_359_123#_c_1489_n 0.00197321f $X=5.3 $Y=2.205
+ $X2=0 $Y2=0
cc_670 N_A_850_51#_c_785_n N_A_359_123#_c_1489_n 0.0522124f $X=4.61 $Y=1.375
+ $X2=0 $Y2=0
cc_671 N_A_850_51#_c_787_n N_A_359_123#_c_1489_n 0.00916142f $X=4.655 $Y=1.4
+ $X2=0 $Y2=0
cc_672 N_A_850_51#_c_795_n N_A_359_123#_c_1489_n 0.0139562f $X=4.61 $Y=1.235
+ $X2=0 $Y2=0
cc_673 N_A_850_51#_c_790_n N_VGND_M1012_d 0.0175919f $X=6.765 $Y=0.64 $X2=0
+ $Y2=0
cc_674 N_A_850_51#_c_796_n N_VGND_M1012_d 0.0104282f $X=6.85 $Y=0.34 $X2=0 $Y2=0
cc_675 N_A_850_51#_c_795_n N_VGND_c_1659_n 8.65947e-19 $X=4.61 $Y=1.235 $X2=0
+ $Y2=0
cc_676 N_A_850_51#_c_788_n N_VGND_c_1672_n 0.0114338f $X=5.72 $Y=0.375 $X2=0
+ $Y2=0
cc_677 N_A_850_51#_c_789_n N_VGND_c_1672_n 0.00648855f $X=5.64 $Y=0.35 $X2=0
+ $Y2=0
cc_678 N_A_850_51#_c_790_n N_VGND_c_1672_n 0.00766817f $X=6.765 $Y=0.64 $X2=0
+ $Y2=0
cc_679 N_A_850_51#_c_794_n N_VGND_c_1672_n 0.0932303f $X=4.665 $Y=0.425 $X2=0
+ $Y2=0
cc_680 N_A_850_51#_c_790_n N_VGND_c_1673_n 0.00378639f $X=6.765 $Y=0.64 $X2=0
+ $Y2=0
cc_681 N_A_850_51#_c_791_n N_VGND_c_1673_n 0.0557663f $X=7.615 $Y=0.34 $X2=0
+ $Y2=0
cc_682 N_A_850_51#_c_796_n N_VGND_c_1673_n 0.0117148f $X=6.85 $Y=0.34 $X2=0
+ $Y2=0
cc_683 N_A_850_51#_c_797_n N_VGND_c_1673_n 0.00313891f $X=7.705 $Y=0.835 $X2=0
+ $Y2=0
cc_684 N_A_850_51#_c_788_n N_VGND_c_1677_n 0.00607686f $X=5.72 $Y=0.375 $X2=0
+ $Y2=0
cc_685 N_A_850_51#_c_789_n N_VGND_c_1677_n 0.00210732f $X=5.64 $Y=0.35 $X2=0
+ $Y2=0
cc_686 N_A_850_51#_c_790_n N_VGND_c_1677_n 0.0243781f $X=6.765 $Y=0.64 $X2=0
+ $Y2=0
cc_687 N_A_850_51#_c_796_n N_VGND_c_1677_n 0.00966701f $X=6.85 $Y=0.34 $X2=0
+ $Y2=0
cc_688 N_A_850_51#_c_788_n N_VGND_c_1680_n 0.00608593f $X=5.72 $Y=0.375 $X2=0
+ $Y2=0
cc_689 N_A_850_51#_c_789_n N_VGND_c_1680_n 0.0100928f $X=5.64 $Y=0.35 $X2=0
+ $Y2=0
cc_690 N_A_850_51#_c_790_n N_VGND_c_1680_n 0.0182197f $X=6.765 $Y=0.64 $X2=0
+ $Y2=0
cc_691 N_A_850_51#_c_791_n N_VGND_c_1680_n 0.0311941f $X=7.615 $Y=0.34 $X2=0
+ $Y2=0
cc_692 N_A_850_51#_c_793_n N_VGND_c_1680_n 0.00197611f $X=7.71 $Y=1 $X2=0 $Y2=0
cc_693 N_A_850_51#_c_794_n N_VGND_c_1680_n 0.0529714f $X=4.665 $Y=0.425 $X2=0
+ $Y2=0
cc_694 N_A_850_51#_c_796_n N_VGND_c_1680_n 0.00646994f $X=6.85 $Y=0.34 $X2=0
+ $Y2=0
cc_695 N_A_850_51#_c_797_n N_VGND_c_1680_n 0.00505852f $X=7.705 $Y=0.835 $X2=0
+ $Y2=0
cc_696 N_A_850_51#_c_788_n A_1143_125# 0.00209416f $X=5.72 $Y=0.375 $X2=-0.19
+ $Y2=-0.245
cc_697 N_A_850_51#_c_790_n A_1143_125# 0.0012269f $X=6.765 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_698 N_A_1203_99#_c_956_n N_A_1053_125#_M1002_g 0.0378647f $X=6.38 $Y=1.58
+ $X2=0 $Y2=0
cc_699 N_A_1203_99#_M1021_g N_A_1053_125#_M1002_g 0.0207383f $X=6.28 $Y=2.455
+ $X2=0 $Y2=0
cc_700 N_A_1203_99#_c_958_n N_A_1053_125#_M1002_g 0.038587f $X=6.92 $Y=1.775
+ $X2=0 $Y2=0
cc_701 N_A_1203_99#_c_960_n N_A_1053_125#_M1002_g 0.00256945f $X=7.36 $Y=1.475
+ $X2=0 $Y2=0
cc_702 N_A_1203_99#_c_960_n N_A_1053_125#_c_1022_n 0.00818835f $X=7.36 $Y=1.475
+ $X2=0 $Y2=0
cc_703 N_A_1203_99#_c_961_n N_A_1053_125#_c_1022_n 0.00922197f $X=7.28 $Y=0.72
+ $X2=0 $Y2=0
cc_704 N_A_1203_99#_c_955_n N_A_1053_125#_c_1023_n 0.00748543f $X=6.09 $Y=1.155
+ $X2=0 $Y2=0
cc_705 N_A_1203_99#_c_956_n N_A_1053_125#_c_1023_n 0.0281811f $X=6.38 $Y=1.58
+ $X2=0 $Y2=0
cc_706 N_A_1203_99#_c_958_n N_A_1053_125#_c_1023_n 0.070168f $X=6.92 $Y=1.775
+ $X2=0 $Y2=0
cc_707 N_A_1203_99#_c_959_n N_A_1053_125#_c_1023_n 3.31618e-19 $X=7.275 $Y=1.565
+ $X2=0 $Y2=0
cc_708 N_A_1203_99#_c_960_n N_A_1053_125#_c_1023_n 0.0189746f $X=7.36 $Y=1.475
+ $X2=0 $Y2=0
cc_709 N_A_1203_99#_c_956_n N_A_1053_125#_c_1025_n 0.00462867f $X=6.38 $Y=1.58
+ $X2=0 $Y2=0
cc_710 N_A_1203_99#_c_955_n N_A_1053_125#_c_1026_n 0.00136843f $X=6.09 $Y=1.155
+ $X2=0 $Y2=0
cc_711 N_A_1203_99#_c_956_n N_A_1053_125#_c_1026_n 0.00713674f $X=6.38 $Y=1.58
+ $X2=0 $Y2=0
cc_712 N_A_1203_99#_c_958_n N_A_1053_125#_c_1026_n 0.00491872f $X=6.92 $Y=1.775
+ $X2=0 $Y2=0
cc_713 N_A_1203_99#_c_959_n N_A_1053_125#_c_1026_n 0.00191333f $X=7.275 $Y=1.565
+ $X2=0 $Y2=0
cc_714 N_A_1203_99#_M1021_g N_VPWR_c_1344_n 6.65218e-19 $X=6.28 $Y=2.455 $X2=0
+ $Y2=0
cc_715 N_A_1203_99#_M1002_d N_VPWR_c_1329_n 0.00283464f $X=6.945 $Y=2.245 $X2=0
+ $Y2=0
cc_716 N_A_1203_99#_c_955_n N_VGND_c_1672_n 0.00316055f $X=6.09 $Y=1.155 $X2=0
+ $Y2=0
cc_717 N_A_1203_99#_c_955_n N_VGND_c_1680_n 0.00469432f $X=6.09 $Y=1.155 $X2=0
+ $Y2=0
cc_718 N_A_1053_125#_M1002_g N_VPWR_c_1345_n 0.00400062f $X=6.87 $Y=2.665 $X2=0
+ $Y2=0
cc_719 N_A_1053_125#_M1002_g N_VPWR_c_1349_n 0.00659856f $X=6.87 $Y=2.665 $X2=0
+ $Y2=0
cc_720 N_A_1053_125#_M1002_g N_VPWR_c_1329_n 0.00686705f $X=6.87 $Y=2.665 $X2=0
+ $Y2=0
cc_721 N_A_1053_125#_c_1049_n N_A_359_123#_c_1488_n 0.0147043f $X=5.425 $Y=0.83
+ $X2=0 $Y2=0
cc_722 N_A_1053_125#_c_1028_n N_A_359_123#_c_1493_n 0.00177665f $X=5.61 $Y=2.48
+ $X2=0 $Y2=0
cc_723 N_A_1053_125#_c_1028_n N_A_359_123#_c_1494_n 0.0116408f $X=5.61 $Y=2.48
+ $X2=0 $Y2=0
cc_724 N_A_1053_125#_c_1024_n N_A_359_123#_c_1489_n 0.0183457f $X=5.32 $Y=1.055
+ $X2=0 $Y2=0
cc_725 N_A_1053_125#_c_1025_n N_A_359_123#_c_1489_n 0.0610848f $X=5.532 $Y=2.225
+ $X2=0 $Y2=0
cc_726 N_A_1053_125#_c_1022_n N_VGND_c_1673_n 0.00313972f $X=7.065 $Y=1.055
+ $X2=0 $Y2=0
cc_727 N_A_1053_125#_c_1022_n N_VGND_c_1677_n 0.00161217f $X=7.065 $Y=1.055
+ $X2=0 $Y2=0
cc_728 N_A_1053_125#_c_1022_n N_VGND_c_1680_n 0.00549465f $X=7.065 $Y=1.055
+ $X2=0 $Y2=0
cc_729 N_A_1673_409#_M1018_g N_A_1475_449#_M1015_g 0.00246637f $X=8.44 $Y=2.745
+ $X2=0 $Y2=0
cc_730 N_A_1673_409#_M1029_g N_A_1475_449#_M1015_g 0.0218348f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_731 N_A_1673_409#_c_1115_n N_A_1475_449#_M1015_g 0.0184565f $X=9.395 $Y=2.13
+ $X2=0 $Y2=0
cc_732 N_A_1673_409#_c_1116_n N_A_1475_449#_M1015_g 0.00208924f $X=9.49 $Y=2.335
+ $X2=0 $Y2=0
cc_733 N_A_1673_409#_c_1118_n N_A_1475_449#_M1015_g 4.49467e-19 $X=8.61 $Y=2.13
+ $X2=0 $Y2=0
cc_734 N_A_1673_409#_M1029_g N_A_1475_449#_c_1251_n 0.00862981f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_735 N_A_1673_409#_M1029_g N_A_1475_449#_c_1240_n 0.00343735f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_736 N_A_1673_409#_c_1118_n N_A_1475_449#_c_1240_n 0.0241314f $X=8.61 $Y=2.13
+ $X2=0 $Y2=0
cc_737 N_A_1673_409#_c_1120_n N_A_1475_449#_c_1240_n 0.00466115f $X=8.7 $Y=2.21
+ $X2=0 $Y2=0
cc_738 N_A_1673_409#_M1029_g N_A_1475_449#_c_1241_n 0.00788485f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_739 N_A_1673_409#_c_1118_n N_A_1475_449#_c_1241_n 0.014816f $X=8.61 $Y=2.13
+ $X2=0 $Y2=0
cc_740 N_A_1673_409#_c_1120_n N_A_1475_449#_c_1241_n 0.00636824f $X=8.7 $Y=2.21
+ $X2=0 $Y2=0
cc_741 N_A_1673_409#_M1029_g N_A_1475_449#_c_1233_n 0.0105013f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_742 N_A_1673_409#_M1029_g N_A_1475_449#_c_1234_n 0.00566284f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_743 N_A_1673_409#_M1029_g N_A_1475_449#_c_1235_n 0.0122546f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_744 N_A_1673_409#_c_1115_n N_A_1475_449#_c_1235_n 0.0155071f $X=9.395 $Y=2.13
+ $X2=0 $Y2=0
cc_745 N_A_1673_409#_c_1102_n N_A_1475_449#_c_1235_n 0.00800193f $X=9.505
+ $Y=1.285 $X2=0 $Y2=0
cc_746 N_A_1673_409#_c_1103_n N_A_1475_449#_c_1235_n 0.0023082f $X=9.49 $Y=1.86
+ $X2=0 $Y2=0
cc_747 N_A_1673_409#_c_1118_n N_A_1475_449#_c_1235_n 0.00114133f $X=8.61 $Y=2.13
+ $X2=0 $Y2=0
cc_748 N_A_1673_409#_c_1106_n N_A_1475_449#_c_1235_n 0.0179024f $X=9.505
+ $Y=1.385 $X2=0 $Y2=0
cc_749 N_A_1673_409#_M1029_g N_A_1475_449#_c_1236_n 0.0213449f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_750 N_A_1673_409#_c_1115_n N_A_1475_449#_c_1236_n 0.00362056f $X=9.395
+ $Y=2.13 $X2=0 $Y2=0
cc_751 N_A_1673_409#_c_1102_n N_A_1475_449#_c_1236_n 0.00122798f $X=9.505
+ $Y=1.285 $X2=0 $Y2=0
cc_752 N_A_1673_409#_c_1103_n N_A_1475_449#_c_1236_n 0.00703443f $X=9.49 $Y=1.86
+ $X2=0 $Y2=0
cc_753 N_A_1673_409#_c_1106_n N_A_1475_449#_c_1236_n 0.00191299f $X=9.505
+ $Y=1.385 $X2=0 $Y2=0
cc_754 N_A_1673_409#_c_1107_n N_A_1475_449#_c_1236_n 0.011868f $X=10.15 $Y=1.37
+ $X2=0 $Y2=0
cc_755 N_A_1673_409#_M1029_g N_A_1475_449#_c_1237_n 0.00653167f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_756 N_A_1673_409#_M1029_g N_A_1475_449#_c_1238_n 0.0167179f $X=8.7 $Y=0.515
+ $X2=0 $Y2=0
cc_757 N_A_1673_409#_c_1102_n N_A_1475_449#_c_1238_n 0.00601686f $X=9.505
+ $Y=1.285 $X2=0 $Y2=0
cc_758 N_A_1673_409#_c_1115_n N_VPWR_M1018_d 0.00695023f $X=9.395 $Y=2.13 $X2=0
+ $Y2=0
cc_759 N_A_1673_409#_M1004_g N_VPWR_c_1333_n 0.00768178f $X=10.225 $Y=2.465
+ $X2=0 $Y2=0
cc_760 N_A_1673_409#_c_1116_n N_VPWR_c_1333_n 0.0450651f $X=9.49 $Y=2.335 $X2=0
+ $Y2=0
cc_761 N_A_1673_409#_c_1103_n N_VPWR_c_1333_n 0.0135605f $X=9.49 $Y=1.86 $X2=0
+ $Y2=0
cc_762 N_A_1673_409#_c_1104_n N_VPWR_c_1333_n 0.0146086f $X=10.85 $Y=1.37 $X2=0
+ $Y2=0
cc_763 N_A_1673_409#_c_1160_p N_VPWR_c_1333_n 0.0110675f $X=9.495 $Y=2.13 $X2=0
+ $Y2=0
cc_764 N_A_1673_409#_c_1107_n N_VPWR_c_1333_n 0.0065947f $X=10.15 $Y=1.37 $X2=0
+ $Y2=0
cc_765 N_A_1673_409#_M1004_g N_VPWR_c_1334_n 7.69681e-19 $X=10.225 $Y=2.465
+ $X2=0 $Y2=0
cc_766 N_A_1673_409#_M1011_g N_VPWR_c_1334_n 0.0163934f $X=10.655 $Y=2.465 $X2=0
+ $Y2=0
cc_767 N_A_1673_409#_M1024_g N_VPWR_c_1334_n 0.0162548f $X=11.085 $Y=2.465 $X2=0
+ $Y2=0
cc_768 N_A_1673_409#_M1036_g N_VPWR_c_1334_n 7.55462e-19 $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_769 N_A_1673_409#_M1024_g N_VPWR_c_1336_n 7.27171e-19 $X=11.085 $Y=2.465
+ $X2=0 $Y2=0
cc_770 N_A_1673_409#_M1036_g N_VPWR_c_1336_n 0.0152814f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_771 N_A_1673_409#_c_1116_n N_VPWR_c_1341_n 0.00866114f $X=9.49 $Y=2.335 $X2=0
+ $Y2=0
cc_772 N_A_1673_409#_M1018_g N_VPWR_c_1345_n 0.00395039f $X=8.44 $Y=2.745 $X2=0
+ $Y2=0
cc_773 N_A_1673_409#_M1004_g N_VPWR_c_1346_n 0.00585385f $X=10.225 $Y=2.465
+ $X2=0 $Y2=0
cc_774 N_A_1673_409#_M1011_g N_VPWR_c_1346_n 0.00486043f $X=10.655 $Y=2.465
+ $X2=0 $Y2=0
cc_775 N_A_1673_409#_M1024_g N_VPWR_c_1347_n 0.00486043f $X=11.085 $Y=2.465
+ $X2=0 $Y2=0
cc_776 N_A_1673_409#_M1036_g N_VPWR_c_1347_n 0.00486043f $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_777 N_A_1673_409#_M1018_g N_VPWR_c_1350_n 0.0116517f $X=8.44 $Y=2.745 $X2=0
+ $Y2=0
cc_778 N_A_1673_409#_c_1115_n N_VPWR_c_1350_n 0.0282638f $X=9.395 $Y=2.13 $X2=0
+ $Y2=0
cc_779 N_A_1673_409#_c_1116_n N_VPWR_c_1350_n 0.0239785f $X=9.49 $Y=2.335 $X2=0
+ $Y2=0
cc_780 N_A_1673_409#_c_1118_n N_VPWR_c_1350_n 0.0140398f $X=8.61 $Y=2.13 $X2=0
+ $Y2=0
cc_781 N_A_1673_409#_c_1120_n N_VPWR_c_1350_n 0.00291024f $X=8.7 $Y=2.21 $X2=0
+ $Y2=0
cc_782 N_A_1673_409#_M1018_g N_VPWR_c_1329_n 0.00471716f $X=8.44 $Y=2.745 $X2=0
+ $Y2=0
cc_783 N_A_1673_409#_M1004_g N_VPWR_c_1329_n 0.0118221f $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_784 N_A_1673_409#_M1011_g N_VPWR_c_1329_n 0.00824727f $X=10.655 $Y=2.465
+ $X2=0 $Y2=0
cc_785 N_A_1673_409#_M1024_g N_VPWR_c_1329_n 0.00824727f $X=11.085 $Y=2.465
+ $X2=0 $Y2=0
cc_786 N_A_1673_409#_M1036_g N_VPWR_c_1329_n 0.00824727f $X=11.515 $Y=2.465
+ $X2=0 $Y2=0
cc_787 N_A_1673_409#_c_1116_n N_VPWR_c_1329_n 0.00729078f $X=9.49 $Y=2.335 $X2=0
+ $Y2=0
cc_788 N_A_1673_409#_M1004_g N_Q_c_1614_n 7.661e-19 $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_789 N_A_1673_409#_M1011_g N_Q_c_1614_n 7.6414e-19 $X=10.655 $Y=2.465 $X2=0
+ $Y2=0
cc_790 N_A_1673_409#_c_1095_n N_Q_c_1605_n 0.0124547f $X=10.655 $Y=1.205 $X2=0
+ $Y2=0
cc_791 N_A_1673_409#_c_1097_n N_Q_c_1605_n 0.0140977f $X=11.085 $Y=1.205 $X2=0
+ $Y2=0
cc_792 N_A_1673_409#_c_1104_n N_Q_c_1605_n 0.0341285f $X=10.85 $Y=1.37 $X2=0
+ $Y2=0
cc_793 N_A_1673_409#_c_1108_n N_Q_c_1605_n 0.00246472f $X=11.515 $Y=1.37 $X2=0
+ $Y2=0
cc_794 N_A_1673_409#_c_1104_n N_Q_c_1606_n 0.0187572f $X=10.85 $Y=1.37 $X2=0
+ $Y2=0
cc_795 N_A_1673_409#_c_1108_n N_Q_c_1606_n 0.00256759f $X=11.515 $Y=1.37 $X2=0
+ $Y2=0
cc_796 N_A_1673_409#_M1011_g N_Q_c_1611_n 0.013997f $X=10.655 $Y=2.465 $X2=0
+ $Y2=0
cc_797 N_A_1673_409#_M1024_g N_Q_c_1611_n 0.0159476f $X=11.085 $Y=2.465 $X2=0
+ $Y2=0
cc_798 N_A_1673_409#_c_1104_n N_Q_c_1611_n 0.0341288f $X=10.85 $Y=1.37 $X2=0
+ $Y2=0
cc_799 N_A_1673_409#_c_1108_n N_Q_c_1611_n 0.00237812f $X=11.515 $Y=1.37 $X2=0
+ $Y2=0
cc_800 N_A_1673_409#_M1004_g N_Q_c_1607_n 0.00544221f $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_801 N_A_1673_409#_c_1104_n N_Q_c_1607_n 0.0183497f $X=10.85 $Y=1.37 $X2=0
+ $Y2=0
cc_802 N_A_1673_409#_c_1108_n N_Q_c_1607_n 0.00247486f $X=11.515 $Y=1.37 $X2=0
+ $Y2=0
cc_803 N_A_1673_409#_c_1099_n N_Q_c_1609_n 0.0129231f $X=11.515 $Y=1.205 $X2=0
+ $Y2=0
cc_804 N_A_1673_409#_M1036_g N_Q_c_1613_n 0.0182711f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_805 N_A_1673_409#_c_1097_n Q 0.00287753f $X=11.085 $Y=1.205 $X2=0 $Y2=0
cc_806 N_A_1673_409#_M1024_g Q 0.00384749f $X=11.085 $Y=2.465 $X2=0 $Y2=0
cc_807 N_A_1673_409#_c_1099_n Q 0.00386991f $X=11.515 $Y=1.205 $X2=0 $Y2=0
cc_808 N_A_1673_409#_M1036_g Q 0.0051892f $X=11.515 $Y=2.465 $X2=0 $Y2=0
cc_809 N_A_1673_409#_c_1104_n Q 0.0159871f $X=10.85 $Y=1.37 $X2=0 $Y2=0
cc_810 N_A_1673_409#_c_1108_n Q 0.0337548f $X=11.515 $Y=1.37 $X2=0 $Y2=0
cc_811 N_A_1673_409#_M1029_g N_VGND_c_1660_n 0.00972994f $X=8.7 $Y=0.515 $X2=0
+ $Y2=0
cc_812 N_A_1673_409#_c_1102_n N_VGND_c_1660_n 5.61173e-19 $X=9.505 $Y=1.285
+ $X2=0 $Y2=0
cc_813 N_A_1673_409#_c_1093_n N_VGND_c_1661_n 0.00702227f $X=10.225 $Y=1.205
+ $X2=0 $Y2=0
cc_814 N_A_1673_409#_c_1101_n N_VGND_c_1661_n 0.0545599f $X=9.44 $Y=0.42 $X2=0
+ $Y2=0
cc_815 N_A_1673_409#_c_1104_n N_VGND_c_1661_n 0.0234825f $X=10.85 $Y=1.37 $X2=0
+ $Y2=0
cc_816 N_A_1673_409#_c_1107_n N_VGND_c_1661_n 0.00739466f $X=10.15 $Y=1.37 $X2=0
+ $Y2=0
cc_817 N_A_1673_409#_c_1093_n N_VGND_c_1662_n 5.8196e-19 $X=10.225 $Y=1.205
+ $X2=0 $Y2=0
cc_818 N_A_1673_409#_c_1095_n N_VGND_c_1662_n 0.0115667f $X=10.655 $Y=1.205
+ $X2=0 $Y2=0
cc_819 N_A_1673_409#_c_1097_n N_VGND_c_1662_n 0.0114291f $X=11.085 $Y=1.205
+ $X2=0 $Y2=0
cc_820 N_A_1673_409#_c_1099_n N_VGND_c_1662_n 5.67983e-19 $X=11.515 $Y=1.205
+ $X2=0 $Y2=0
cc_821 N_A_1673_409#_c_1097_n N_VGND_c_1664_n 5.67983e-19 $X=11.085 $Y=1.205
+ $X2=0 $Y2=0
cc_822 N_A_1673_409#_c_1099_n N_VGND_c_1664_n 0.0140537f $X=11.515 $Y=1.205
+ $X2=0 $Y2=0
cc_823 N_A_1673_409#_c_1101_n N_VGND_c_1669_n 0.0178111f $X=9.44 $Y=0.42 $X2=0
+ $Y2=0
cc_824 N_A_1673_409#_M1029_g N_VGND_c_1673_n 0.00442016f $X=8.7 $Y=0.515 $X2=0
+ $Y2=0
cc_825 N_A_1673_409#_c_1093_n N_VGND_c_1674_n 0.00565115f $X=10.225 $Y=1.205
+ $X2=0 $Y2=0
cc_826 N_A_1673_409#_c_1095_n N_VGND_c_1674_n 0.00469214f $X=10.655 $Y=1.205
+ $X2=0 $Y2=0
cc_827 N_A_1673_409#_c_1097_n N_VGND_c_1675_n 0.00469214f $X=11.085 $Y=1.205
+ $X2=0 $Y2=0
cc_828 N_A_1673_409#_c_1099_n N_VGND_c_1675_n 0.00469214f $X=11.515 $Y=1.205
+ $X2=0 $Y2=0
cc_829 N_A_1673_409#_M1013_d N_VGND_c_1680_n 0.00371702f $X=9.3 $Y=0.235 $X2=0
+ $Y2=0
cc_830 N_A_1673_409#_M1029_g N_VGND_c_1680_n 0.00808394f $X=8.7 $Y=0.515 $X2=0
+ $Y2=0
cc_831 N_A_1673_409#_c_1093_n N_VGND_c_1680_n 0.0117308f $X=10.225 $Y=1.205
+ $X2=0 $Y2=0
cc_832 N_A_1673_409#_c_1095_n N_VGND_c_1680_n 0.00825323f $X=10.655 $Y=1.205
+ $X2=0 $Y2=0
cc_833 N_A_1673_409#_c_1097_n N_VGND_c_1680_n 0.00825323f $X=11.085 $Y=1.205
+ $X2=0 $Y2=0
cc_834 N_A_1673_409#_c_1099_n N_VGND_c_1680_n 0.00825323f $X=11.515 $Y=1.205
+ $X2=0 $Y2=0
cc_835 N_A_1673_409#_c_1101_n N_VGND_c_1680_n 0.0100304f $X=9.44 $Y=0.42 $X2=0
+ $Y2=0
cc_836 N_A_1475_449#_M1015_g N_VPWR_c_1333_n 0.00381281f $X=9.275 $Y=2.325 $X2=0
+ $Y2=0
cc_837 N_A_1475_449#_M1015_g N_VPWR_c_1341_n 0.00379792f $X=9.275 $Y=2.325 $X2=0
+ $Y2=0
cc_838 N_A_1475_449#_c_1247_n N_VPWR_c_1345_n 0.0158342f $X=8.155 $Y=2.745 $X2=0
+ $Y2=0
cc_839 N_A_1475_449#_M1015_g N_VPWR_c_1350_n 0.0119889f $X=9.275 $Y=2.325 $X2=0
+ $Y2=0
cc_840 N_A_1475_449#_c_1240_n N_VPWR_c_1350_n 0.00513665f $X=8.24 $Y=2.58 $X2=0
+ $Y2=0
cc_841 N_A_1475_449#_M1023_d N_VPWR_c_1329_n 0.0033464f $X=7.375 $Y=2.245 $X2=0
+ $Y2=0
cc_842 N_A_1475_449#_M1015_g N_VPWR_c_1329_n 0.00453573f $X=9.275 $Y=2.325 $X2=0
+ $Y2=0
cc_843 N_A_1475_449#_c_1247_n N_VPWR_c_1329_n 0.0184776f $X=8.155 $Y=2.745 $X2=0
+ $Y2=0
cc_844 N_A_1475_449#_c_1247_n A_1631_507# 0.00128978f $X=8.155 $Y=2.745
+ $X2=-0.19 $Y2=-0.245
cc_845 N_A_1475_449#_c_1251_n N_VGND_c_1660_n 0.0272528f $X=8.515 $Y=0.51 $X2=0
+ $Y2=0
cc_846 N_A_1475_449#_c_1233_n N_VGND_c_1660_n 0.0254949f $X=8.6 $Y=1.185 $X2=0
+ $Y2=0
cc_847 N_A_1475_449#_c_1235_n N_VGND_c_1660_n 0.0241758f $X=9.15 $Y=1.35 $X2=0
+ $Y2=0
cc_848 N_A_1475_449#_c_1236_n N_VGND_c_1660_n 0.0036701f $X=9.15 $Y=1.35 $X2=0
+ $Y2=0
cc_849 N_A_1475_449#_c_1238_n N_VGND_c_1660_n 0.0143441f $X=9.167 $Y=1.185 $X2=0
+ $Y2=0
cc_850 N_A_1475_449#_c_1238_n N_VGND_c_1661_n 0.00276642f $X=9.167 $Y=1.185
+ $X2=0 $Y2=0
cc_851 N_A_1475_449#_c_1238_n N_VGND_c_1669_n 0.00486043f $X=9.167 $Y=1.185
+ $X2=0 $Y2=0
cc_852 N_A_1475_449#_c_1251_n N_VGND_c_1673_n 0.0269111f $X=8.515 $Y=0.51 $X2=0
+ $Y2=0
cc_853 N_A_1475_449#_c_1251_n N_VGND_c_1680_n 0.0251663f $X=8.515 $Y=0.51 $X2=0
+ $Y2=0
cc_854 N_A_1475_449#_c_1238_n N_VGND_c_1680_n 0.00954696f $X=9.167 $Y=1.185
+ $X2=0 $Y2=0
cc_855 N_A_1475_449#_c_1251_n A_1670_61# 0.00604812f $X=8.515 $Y=0.51 $X2=-0.19
+ $Y2=-0.245
cc_856 N_A_1475_449#_c_1233_n A_1670_61# 5.66458e-19 $X=8.6 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_857 N_VPWR_c_1329_n A_296_491# 0.00314438f $X=11.76 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_858 N_VPWR_c_1329_n N_A_359_123#_M1020_d 0.00236474f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_859 N_VPWR_c_1330_n N_A_359_123#_c_1497_n 0.0116395f $X=1.19 $Y=2.805 $X2=0
+ $Y2=0
cc_860 N_VPWR_c_1331_n N_A_359_123#_c_1497_n 0.0245556f $X=2.915 $Y=2.825 $X2=0
+ $Y2=0
cc_861 N_VPWR_c_1337_n N_A_359_123#_c_1497_n 0.0288353f $X=2.82 $Y=3.33 $X2=0
+ $Y2=0
cc_862 N_VPWR_c_1329_n N_A_359_123#_c_1497_n 0.0288974f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_863 N_VPWR_M1001_d N_A_359_123#_c_1491_n 0.00167354f $X=2.74 $Y=2.455 $X2=0
+ $Y2=0
cc_864 N_VPWR_M1003_s N_A_359_123#_c_1491_n 0.00826046f $X=3.74 $Y=2.405 $X2=0
+ $Y2=0
cc_865 N_VPWR_c_1331_n N_A_359_123#_c_1491_n 0.00157285f $X=2.915 $Y=2.825 $X2=0
+ $Y2=0
cc_866 N_VPWR_c_1332_n N_A_359_123#_c_1491_n 0.00678346f $X=3.865 $Y=2.805 $X2=0
+ $Y2=0
cc_867 N_VPWR_M1001_d N_A_359_123#_c_1502_n 0.00214811f $X=2.74 $Y=2.455 $X2=0
+ $Y2=0
cc_868 N_VPWR_M1001_d N_A_359_123#_c_1492_n 0.00243619f $X=2.74 $Y=2.455 $X2=0
+ $Y2=0
cc_869 N_VPWR_c_1331_n N_A_359_123#_c_1492_n 0.0137758f $X=2.915 $Y=2.825 $X2=0
+ $Y2=0
cc_870 N_VPWR_c_1329_n N_A_359_123#_c_1492_n 0.00502602f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_871 N_VPWR_c_1329_n A_454_491# 0.00270181f $X=11.76 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_872 N_VPWR_c_1329_n N_Q_M1004_s 0.0041489f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_873 N_VPWR_c_1329_n N_Q_M1024_s 0.00536646f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_874 N_VPWR_c_1333_n N_Q_c_1614_n 6.8221e-19 $X=10.01 $Y=1.98 $X2=0 $Y2=0
cc_875 N_VPWR_c_1346_n N_Q_c_1614_n 0.0136943f $X=10.705 $Y=3.33 $X2=0 $Y2=0
cc_876 N_VPWR_c_1329_n N_Q_c_1614_n 0.00866972f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_877 N_VPWR_c_1334_n N_Q_c_1611_n 0.0216087f $X=10.87 $Y=2.08 $X2=0 $Y2=0
cc_878 N_VPWR_c_1333_n N_Q_c_1607_n 8.76939e-19 $X=10.01 $Y=1.98 $X2=0 $Y2=0
cc_879 N_VPWR_c_1347_n N_Q_c_1644_n 0.0124525f $X=11.565 $Y=3.33 $X2=0 $Y2=0
cc_880 N_VPWR_c_1329_n N_Q_c_1644_n 0.00730901f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_881 N_VPWR_M1036_d N_Q_c_1613_n 0.00272521f $X=11.59 $Y=1.835 $X2=0 $Y2=0
cc_882 N_VPWR_c_1336_n N_Q_c_1613_n 0.0243971f $X=11.73 $Y=2.18 $X2=0 $Y2=0
cc_883 N_A_359_123#_c_1497_n A_454_491# 0.00730063f $X=2.48 $Y=2.805 $X2=-0.19
+ $Y2=-0.245
cc_884 N_A_359_123#_c_1500_n A_454_491# 0.0017662f $X=2.565 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_885 N_A_359_123#_c_1492_n A_454_491# 3.96176e-19 $X=2.64 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_886 N_A_359_123#_c_1508_n N_VGND_c_1658_n 0.00403364f $X=2.03 $Y=0.89 $X2=0
+ $Y2=0
cc_887 N_A_359_123#_c_1485_n N_VGND_c_1658_n 0.0228102f $X=2.905 $Y=1.13 $X2=0
+ $Y2=0
cc_888 N_A_359_123#_c_1508_n N_VGND_c_1667_n 0.00293619f $X=2.03 $Y=0.89 $X2=0
+ $Y2=0
cc_889 N_A_359_123#_c_1508_n N_VGND_c_1680_n 0.00452458f $X=2.03 $Y=0.89 $X2=0
+ $Y2=0
cc_890 N_Q_c_1605_n N_VGND_M1014_d 0.00176461f $X=11.195 $Y=1.03 $X2=0 $Y2=0
cc_891 N_Q_c_1609_n N_VGND_M1025_d 0.00300749f $X=11.552 $Y=1.03 $X2=0 $Y2=0
cc_892 N_Q_c_1606_n N_VGND_c_1661_n 0.00166417f $X=10.535 $Y=1.03 $X2=0 $Y2=0
cc_893 N_Q_c_1605_n N_VGND_c_1662_n 0.0170777f $X=11.195 $Y=1.03 $X2=0 $Y2=0
cc_894 N_Q_c_1609_n N_VGND_c_1664_n 0.0243971f $X=11.552 $Y=1.03 $X2=0 $Y2=0
cc_895 N_Q_c_1604_n N_VGND_c_1674_n 0.0138717f $X=10.44 $Y=0.42 $X2=0 $Y2=0
cc_896 N_Q_c_1608_n N_VGND_c_1675_n 0.0124525f $X=11.3 $Y=0.42 $X2=0 $Y2=0
cc_897 N_Q_c_1604_n N_VGND_c_1680_n 0.00886411f $X=10.44 $Y=0.42 $X2=0 $Y2=0
cc_898 N_Q_c_1608_n N_VGND_c_1680_n 0.00730901f $X=11.3 $Y=0.42 $X2=0 $Y2=0
