* File: sky130_fd_sc_lp__a41oi_0.pex.spice
* Created: Wed Sep  2 09:29:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41OI_0%B1 3 6 9 13 15 16 20
r37 20 23 87.7315 $w=4.7e-07 $l=5.05e-07 $layer=POLY_cond $X=0.405 $Y=0.99
+ $X2=0.405 $Y2=1.495
r38 20 22 47.4991 $w=4.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=0.99
+ $X2=0.405 $Y2=0.825
r39 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.335
+ $Y=0.99 $X2=0.335 $Y2=0.99
r40 16 21 9.63 $w=3.63e-07 $l=3.05e-07 $layer=LI1_cond $X=0.267 $Y=1.295
+ $X2=0.267 $Y2=0.99
r41 15 21 2.0523 $w=3.63e-07 $l=6.5e-08 $layer=LI1_cond $X=0.267 $Y=0.925
+ $X2=0.267 $Y2=0.99
r42 11 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.565 $Y=1.81
+ $X2=0.805 $Y2=1.81
r43 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.805 $Y=1.885
+ $X2=0.805 $Y2=1.81
r44 7 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=0.805 $Y=1.885
+ $X2=0.805 $Y2=2.715
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=1.735
+ $X2=0.565 $Y2=1.81
r46 6 23 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.565 $Y=1.735
+ $X2=0.565 $Y2=1.495
r47 3 22 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.565 $Y=0.445
+ $X2=0.565 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%A1 2 5 11 13 14 15 16 17 18 23
c49 15 0 3.2985e-19 $X=1.2 $Y=1.885
r50 23 25 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=0.99
+ $X2=1.06 $Y2=0.825
r51 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.075
+ $Y=0.99 $X2=1.075 $Y2=0.99
r52 17 18 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.295
+ $X2=1.175 $Y2=1.665
r53 17 24 9.49987 $w=3.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.175 $Y=1.295
+ $X2=1.175 $Y2=0.99
r54 16 24 2.02456 $w=3.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.175 $Y=0.925
+ $X2=1.175 $Y2=0.99
r55 14 15 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.2 $Y=1.735 $X2=1.2
+ $Y2=1.885
r56 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.165 $Y=1.495
+ $X2=1.165 $Y2=1.735
r57 11 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.235 $Y=2.715
+ $X2=1.235 $Y2=1.885
r58 5 25 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.075 $Y=0.445
+ $X2=1.075 $Y2=0.825
r59 2 13 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.06 $Y=1.315 $X2=1.06
+ $Y2=1.495
r60 1 23 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.06 $Y=1.005
+ $X2=1.06 $Y2=0.99
r61 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.06 $Y=1.005 $X2=1.06
+ $Y2=1.315
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%A2 3 7 11 12 13 14 15 20
c42 12 0 1.33876e-19 $X=1.615 $Y=1.495
r43 14 15 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.692 $Y=1.295
+ $X2=1.692 $Y2=1.665
r44 13 14 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.692 $Y=0.925
+ $X2=1.692 $Y2=1.295
r45 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.615
+ $Y=0.99 $X2=1.615 $Y2=0.99
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.615 $Y=1.33
+ $X2=1.615 $Y2=0.99
r47 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.33
+ $X2=1.615 $Y2=1.495
r48 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=0.825
+ $X2=1.615 $Y2=0.99
r49 7 12 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=1.665 $Y=2.715
+ $X2=1.665 $Y2=1.495
r50 3 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.525 $Y=0.445
+ $X2=1.525 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%A3 3 7 11 12 13 14 15 20
r42 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=1.295
+ $X2=2.19 $Y2=1.665
r43 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=0.925
+ $X2=2.19 $Y2=1.295
r44 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.185
+ $Y=0.99 $X2=2.185 $Y2=0.99
r45 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.185 $Y=1.33
+ $X2=2.185 $Y2=0.99
r46 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.185 $Y=1.33
+ $X2=2.185 $Y2=1.495
r47 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.185 $Y=0.825
+ $X2=2.185 $Y2=0.99
r48 7 12 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.095 $Y=2.715
+ $X2=2.095 $Y2=1.495
r49 3 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.095 $Y=0.445
+ $X2=2.095 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%A4 3 7 10 13 17 18 19 21 28
r36 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.755
+ $Y=1.08 $X2=2.755 $Y2=1.08
r37 21 29 5.16649 $w=8.43e-07 $l=3.65e-07 $layer=LI1_cond $X=3.12 $Y=1.417
+ $X2=2.755 $Y2=1.417
r38 19 29 1.6278 $w=8.43e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.417
+ $X2=2.755 $Y2=1.417
r39 17 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.755 $Y=1.42
+ $X2=2.755 $Y2=1.08
r40 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.42
+ $X2=2.755 $Y2=1.585
r41 16 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=0.915
+ $X2=2.755 $Y2=1.08
r42 11 13 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.525 $Y=1.81
+ $X2=2.665 $Y2=1.81
r43 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.665 $Y=1.735
+ $X2=2.665 $Y2=1.81
r44 10 18 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.665 $Y=1.735
+ $X2=2.665 $Y2=1.585
r45 7 16 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.665 $Y=0.445 $X2=2.665
+ $Y2=0.915
r46 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.525 $Y=1.885
+ $X2=2.525 $Y2=1.81
r47 1 3 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.525 $Y=1.885
+ $X2=2.525 $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%Y 1 2 9 11 13 14 15 16 17 18
c41 14 0 1.87411e-19 $X=0.622 $Y=1.855
c42 13 0 1.83885e-19 $X=0.622 $Y=1.685
c43 9 0 1.42439e-19 $X=0.59 $Y=2.54
r44 17 18 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.467
+ $X2=2.16 $Y2=0.467
r45 16 17 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.467
+ $X2=1.68 $Y2=0.467
r46 16 23 11.6781 $w=3.73e-07 $l=3.8e-07 $layer=LI1_cond $X=1.2 $Y=0.467
+ $X2=0.82 $Y2=0.467
r47 15 23 2.66378 $w=3.75e-07 $l=1e-07 $layer=LI1_cond $X=0.72 $Y=0.467 $X2=0.82
+ $Y2=0.467
r48 13 14 7.84278 $w=2.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.622 $Y=1.685
+ $X2=0.622 $Y2=1.855
r49 11 15 5.0079 $w=2e-07 $l=1.88e-07 $layer=LI1_cond $X=0.72 $Y=0.655 $X2=0.72
+ $Y2=0.467
r50 11 13 57.1182 $w=1.98e-07 $l=1.03e-06 $layer=LI1_cond $X=0.72 $Y=0.655
+ $X2=0.72 $Y2=1.685
r51 9 14 26.7601 $w=2.93e-07 $l=6.85e-07 $layer=LI1_cond $X=0.572 $Y=2.54
+ $X2=0.572 $Y2=1.855
r52 2 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.465
+ $Y=2.395 $X2=0.59 $Y2=2.54
r53 1 15 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.235 $X2=0.8 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%A_176_479# 1 2 3 12 14 15 18 20 24 26
c44 26 0 1.33876e-19 $X=1.875 $Y=2.115
r45 22 24 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.76 $Y=2.205
+ $X2=2.76 $Y2=2.54
r46 21 26 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=2.005 $Y=2.115
+ $X2=1.875 $Y2=2.115
r47 20 22 7.31368 $w=1.8e-07 $l=1.84594e-07 $layer=LI1_cond $X=2.615 $Y=2.115
+ $X2=2.76 $Y2=2.205
r48 20 21 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=2.615 $Y=2.115
+ $X2=2.005 $Y2=2.115
r49 16 26 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=1.875 $Y=2.205
+ $X2=1.875 $Y2=2.115
r50 16 18 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.875 $Y=2.205
+ $X2=1.875 $Y2=2.54
r51 14 26 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=1.745 $Y=2.115
+ $X2=1.875 $Y2=2.115
r52 14 15 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=1.745 $Y=2.115
+ $X2=1.15 $Y2=2.115
r53 10 15 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=1.02 $Y=2.205
+ $X2=1.15 $Y2=2.115
r54 10 12 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.02 $Y=2.205
+ $X2=1.02 $Y2=2.54
r55 3 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.6
+ $Y=2.395 $X2=2.74 $Y2=2.54
r56 2 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.74
+ $Y=2.395 $X2=1.88 $Y2=2.54
r57 1 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.88
+ $Y=2.395 $X2=1.02 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%VPWR 1 2 9 13 16 17 19 20 21 34 35
r37 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 19 31 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 19 20 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.31 $Y2=3.33
r48 18 34 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 18 20 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.31 $Y2=3.33
r50 16 28 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.32 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 16 17 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.447 $Y2=3.33
r52 15 31 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 15 17 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.447 $Y2=3.33
r54 11 20 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=3.245
+ $X2=2.31 $Y2=3.33
r55 11 13 30.0916 $w=2.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.31 $Y=3.245
+ $X2=2.31 $Y2=2.54
r56 7 17 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.447 $Y=3.245
+ $X2=1.447 $Y2=3.33
r57 7 9 31.8617 $w=2.53e-07 $l=7.05e-07 $layer=LI1_cond $X=1.447 $Y=3.245
+ $X2=1.447 $Y2=2.54
r58 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.17
+ $Y=2.395 $X2=2.31 $Y2=2.54
r59 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.31
+ $Y=2.395 $X2=1.45 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_0%VGND 1 2 7 9 13 16 17 18 28 29
r35 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 26 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r38 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r40 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r41 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 20 32 3.59063 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.225
+ $Y2=0
r43 20 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.72
+ $Y2=0
r44 18 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r45 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r46 16 25 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.64
+ $Y2=0
r47 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.88
+ $Y2=0
r48 15 28 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.12
+ $Y2=0
r49 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=2.88
+ $Y2=0
r50 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0
r51 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0.445
r52 7 32 3.30338 $w=2.05e-07 $l=1.58915e-07 $layer=LI1_cond $X=0.347 $Y=0.085
+ $X2=0.225 $Y2=0
r53 7 9 19.4767 $w=2.03e-07 $l=3.6e-07 $layer=LI1_cond $X=0.347 $Y=0.085
+ $X2=0.347 $Y2=0.445
r54 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.74
+ $Y=0.235 $X2=2.88 $Y2=0.445
r55 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.235 $X2=0.35 $Y2=0.445
.ends

