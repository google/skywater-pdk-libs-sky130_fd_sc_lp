* File: sky130_fd_sc_lp__nor3_1.pxi.spice
* Created: Fri Aug 28 10:55:19 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3_1%A N_A_M1002_g N_A_M1005_g A A N_A_c_40_n N_A_c_41_n
+ PM_SKY130_FD_SC_LP__NOR3_1%A
x_PM_SKY130_FD_SC_LP__NOR3_1%B N_B_M1003_g N_B_M1004_g B B B B N_B_c_64_n
+ N_B_c_65_n B PM_SKY130_FD_SC_LP__NOR3_1%B
x_PM_SKY130_FD_SC_LP__NOR3_1%C N_C_M1001_g N_C_M1000_g C N_C_c_109_n
+ PM_SKY130_FD_SC_LP__NOR3_1%C
x_PM_SKY130_FD_SC_LP__NOR3_1%VPWR N_VPWR_M1005_s N_VPWR_c_135_n N_VPWR_c_136_n
+ VPWR N_VPWR_c_137_n N_VPWR_c_134_n VPWR PM_SKY130_FD_SC_LP__NOR3_1%VPWR
x_PM_SKY130_FD_SC_LP__NOR3_1%Y N_Y_M1002_d N_Y_M1001_d N_Y_M1000_d N_Y_c_202_p
+ N_Y_c_168_n N_Y_c_171_n N_Y_c_162_n N_Y_c_163_n N_Y_c_164_n Y Y Y
+ PM_SKY130_FD_SC_LP__NOR3_1%Y
x_PM_SKY130_FD_SC_LP__NOR3_1%VGND N_VGND_M1002_s N_VGND_M1003_d N_VGND_c_208_n
+ N_VGND_c_209_n N_VGND_c_210_n VGND N_VGND_c_211_n N_VGND_c_212_n
+ N_VGND_c_213_n N_VGND_c_214_n VGND PM_SKY130_FD_SC_LP__NOR3_1%VGND
cc_1 VNB N_A_M1005_g 0.00692274f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB A 0.0200523f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_40_n 0.0385413f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_4 VNB N_A_c_41_n 0.022684f $X=-0.19 $Y=-0.245 $X2=0.377 $Y2=1.21
cc_5 VNB N_B_M1003_g 0.0250691f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.665
cc_6 VNB N_B_c_64_n 0.0240848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_65_n 0.00456739f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_8 VNB N_C_M1001_g 0.0300334f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.665
cc_9 VNB C 0.0225282f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_C_c_109_n 0.0364397f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_11 VNB N_VPWR_c_134_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_Y_c_162_n 0.00435796f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_Y_c_163_n 0.00745959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_164_n 0.0237221f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_15 VNB N_VGND_c_208_n 0.0104415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_209_n 0.0341436f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_VGND_c_210_n 6.14598e-19 $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_18 VNB N_VGND_c_211_n 0.0135197f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_19 VNB N_VGND_c_212_n 0.0181175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_213_n 0.130856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_214_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A_M1005_g 0.0257409f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_23 VPB A 0.00697301f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_24 VPB N_B_M1004_g 0.0187857f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB B 0.00123015f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_26 VPB N_B_c_64_n 0.00817499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_C_M1000_g 0.0255466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB C 0.00366132f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_29 VPB N_C_c_109_n 0.0106067f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_30 VPB N_VPWR_c_135_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.54
cc_31 VPB N_VPWR_c_136_n 0.0484529f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_32 VPB N_VPWR_c_137_n 0.042755f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_33 VPB N_VPWR_c_134_n 0.0441318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_Y_c_162_n 0.00123753f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_35 VPB Y 0.0155303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB Y 0.0400072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 A N_B_M1003_g 6.9343e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_38 N_A_c_41_n N_B_M1003_g 0.0215005f $X=0.377 $Y=1.21 $X2=0 $Y2=0
cc_39 N_A_M1005_g N_B_M1004_g 0.0564527f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_40 N_A_M1005_g B 0.00755325f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_41 A N_B_c_64_n 2.74217e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_42 N_A_c_40_n N_B_c_64_n 0.0199673f $X=0.37 $Y=1.375 $X2=0 $Y2=0
cc_43 A N_B_c_65_n 0.0324943f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_44 N_A_c_40_n N_B_c_65_n 0.00755325f $X=0.37 $Y=1.375 $X2=0 $Y2=0
cc_45 N_A_M1005_g N_VPWR_c_136_n 0.0236354f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_46 A N_VPWR_c_136_n 0.026915f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A_c_40_n N_VPWR_c_136_n 8.38351e-19 $X=0.37 $Y=1.375 $X2=0 $Y2=0
cc_48 N_A_M1005_g N_VPWR_c_137_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_49 N_A_M1005_g N_VPWR_c_134_n 0.00845871f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_50 A N_VGND_c_209_n 0.0260595f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A_c_40_n N_VGND_c_209_n 0.00137064f $X=0.37 $Y=1.375 $X2=0 $Y2=0
cc_52 N_A_c_41_n N_VGND_c_209_n 0.0164545f $X=0.377 $Y=1.21 $X2=0 $Y2=0
cc_53 N_A_c_41_n N_VGND_c_210_n 5.3764e-19 $X=0.377 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A_c_41_n N_VGND_c_211_n 0.00477554f $X=0.377 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A_c_41_n N_VGND_c_213_n 0.00828349f $X=0.377 $Y=1.21 $X2=0 $Y2=0
cc_56 N_B_M1003_g N_C_M1001_g 0.0303755f $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_57 N_B_M1004_g N_C_M1000_g 0.0621559f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_58 B N_C_M1000_g 0.002786f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_59 N_B_c_64_n N_C_c_109_n 0.0204656f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_60 N_B_c_65_n N_C_c_109_n 2.90565e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_61 N_B_M1004_g N_VPWR_c_136_n 0.00257581f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_62 B N_VPWR_c_136_n 0.067972f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_63 N_B_M1004_g N_VPWR_c_137_n 0.00527211f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_64 B N_VPWR_c_137_n 0.00883036f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_65 N_B_M1004_g N_VPWR_c_134_n 0.00954407f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_66 B N_VPWR_c_134_n 0.00970302f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_67 B A_110_367# 0.0153451f $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_68 N_B_M1003_g N_Y_c_168_n 0.0136751f $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_69 N_B_c_64_n N_Y_c_168_n 0.00221742f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_70 N_B_c_65_n N_Y_c_168_n 0.00826538f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_71 N_B_c_64_n N_Y_c_171_n 2.03309e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_72 N_B_c_65_n N_Y_c_171_n 0.00965377f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_73 N_B_M1003_g N_Y_c_162_n 0.00619906f $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_74 N_B_M1004_g N_Y_c_162_n 0.00115341f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_75 B N_Y_c_162_n 0.00851274f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_76 N_B_c_64_n N_Y_c_162_n 0.00204642f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_77 N_B_c_65_n N_Y_c_162_n 0.0254366f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_78 N_B_M1004_g Y 0.00256834f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_79 B Y 0.0178882f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_80 N_B_M1004_g Y 0.00295974f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_81 B Y 0.0229578f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_82 N_B_M1003_g N_VGND_c_209_n 6.13753e-19 $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_83 N_B_M1003_g N_VGND_c_210_n 0.00899708f $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_84 N_B_M1003_g N_VGND_c_211_n 0.00554242f $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_85 N_B_M1003_g N_VGND_c_213_n 0.0095208f $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_86 N_C_M1000_g N_VPWR_c_137_n 0.0054895f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_87 N_C_M1000_g N_VPWR_c_134_n 0.0110663f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_88 N_C_M1001_g N_Y_c_162_n 0.0113042f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_89 N_C_M1000_g N_Y_c_162_n 0.00845186f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_90 C N_Y_c_162_n 0.0335971f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_91 N_C_c_109_n N_Y_c_162_n 0.0076458f $X=1.605 $Y=1.51 $X2=0 $Y2=0
cc_92 N_C_M1001_g N_Y_c_163_n 0.0155203f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_93 C N_Y_c_163_n 0.0188989f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_94 N_C_c_109_n N_Y_c_163_n 0.00263177f $X=1.605 $Y=1.51 $X2=0 $Y2=0
cc_95 N_C_M1000_g Y 0.0176318f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_96 C Y 0.0254492f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_C_c_109_n Y 0.00355733f $X=1.605 $Y=1.51 $X2=0 $Y2=0
cc_98 N_C_M1000_g Y 0.0194747f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_99 N_C_M1001_g N_VGND_c_210_n 0.0105353f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_100 N_C_M1001_g N_VGND_c_212_n 0.00554242f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_101 N_C_M1001_g N_VGND_c_213_n 0.0104879f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_102 N_VPWR_c_134_n A_110_367# 0.00531213f $X=1.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_103 N_VPWR_c_134_n A_202_367# 0.0124205f $X=1.68 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_104 N_VPWR_c_134_n N_Y_M1000_d 0.00215158f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_105 N_VPWR_c_137_n Y 0.0267816f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_106 N_VPWR_c_134_n Y 0.0156791f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_107 A_202_367# N_Y_c_162_n 2.84889e-19 $X=1.01 $Y=1.835 $X2=1.68 $Y2=3.33
cc_108 A_202_367# Y 0.00610199f $X=1.01 $Y=1.835 $X2=0.72 $Y2=3.33
cc_109 N_Y_c_168_n N_VGND_M1003_d 0.00558993f $X=1.18 $Y=0.955 $X2=0 $Y2=0
cc_110 N_Y_c_162_n N_VGND_M1003_d 7.16347e-19 $X=1.265 $Y=1.845 $X2=0 $Y2=0
cc_111 N_Y_c_163_n N_VGND_M1003_d 8.5303e-19 $X=1.615 $Y=0.87 $X2=0 $Y2=0
cc_112 N_Y_c_168_n N_VGND_c_210_n 0.0172485f $X=1.18 $Y=0.955 $X2=0 $Y2=0
cc_113 N_Y_c_202_p N_VGND_c_211_n 0.0131621f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_114 N_Y_c_164_n N_VGND_c_212_n 0.0183924f $X=1.59 $Y=0.42 $X2=0 $Y2=0
cc_115 N_Y_M1002_d N_VGND_c_213_n 0.00467071f $X=0.55 $Y=0.245 $X2=0 $Y2=0
cc_116 N_Y_M1001_d N_VGND_c_213_n 0.00299269f $X=1.45 $Y=0.245 $X2=0 $Y2=0
cc_117 N_Y_c_202_p N_VGND_c_213_n 0.00808656f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_118 N_Y_c_164_n N_VGND_c_213_n 0.0107796f $X=1.59 $Y=0.42 $X2=0 $Y2=0
