* File: sky130_fd_sc_lp__o22a_4.pxi.spice
* Created: Fri Aug 28 11:09:53 2020
* 
x_PM_SKY130_FD_SC_LP__O22A_4%A_86_23# N_A_86_23#_M1010_d N_A_86_23#_M1021_d
+ N_A_86_23#_M1008_s N_A_86_23#_M1001_d N_A_86_23#_M1005_g N_A_86_23#_M1011_g
+ N_A_86_23#_M1002_g N_A_86_23#_M1015_g N_A_86_23#_M1009_g N_A_86_23#_M1016_g
+ N_A_86_23#_M1014_g N_A_86_23#_M1022_g N_A_86_23#_c_180_p N_A_86_23#_c_102_n
+ N_A_86_23#_c_103_n N_A_86_23#_c_104_n N_A_86_23#_c_105_n N_A_86_23#_c_115_p
+ N_A_86_23#_c_157_p N_A_86_23#_c_119_p N_A_86_23#_c_106_n N_A_86_23#_c_117_p
+ N_A_86_23#_c_146_p N_A_86_23#_c_107_n PM_SKY130_FD_SC_LP__O22A_4%A_86_23#
x_PM_SKY130_FD_SC_LP__O22A_4%B1 N_B1_M1010_g N_B1_M1003_g N_B1_M1019_g
+ N_B1_M1023_g N_B1_c_248_n N_B1_c_249_n N_B1_c_250_n N_B1_c_251_n B1
+ N_B1_c_252_n N_B1_c_253_n N_B1_c_254_n PM_SKY130_FD_SC_LP__O22A_4%B1
x_PM_SKY130_FD_SC_LP__O22A_4%B2 N_B2_M1006_g N_B2_M1008_g N_B2_M1021_g
+ N_B2_M1018_g B2 N_B2_c_332_n N_B2_c_329_n PM_SKY130_FD_SC_LP__O22A_4%B2
x_PM_SKY130_FD_SC_LP__O22A_4%A1 N_A1_M1000_g N_A1_M1007_g N_A1_M1012_g
+ N_A1_M1013_g N_A1_c_374_n N_A1_c_375_n N_A1_c_376_n A1 A1 N_A1_c_378_n
+ N_A1_c_379_n N_A1_c_380_n PM_SKY130_FD_SC_LP__O22A_4%A1
x_PM_SKY130_FD_SC_LP__O22A_4%A2 N_A2_M1004_g N_A2_M1001_g N_A2_M1020_g
+ N_A2_M1017_g A2 N_A2_c_446_n PM_SKY130_FD_SC_LP__O22A_4%A2
x_PM_SKY130_FD_SC_LP__O22A_4%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_M1022_d
+ N_VPWR_M1023_s N_VPWR_M1013_d N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n
+ N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n
+ N_VPWR_c_499_n VPWR N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_490_n
+ PM_SKY130_FD_SC_LP__O22A_4%VPWR
x_PM_SKY130_FD_SC_LP__O22A_4%X N_X_M1005_d N_X_M1015_d N_X_M1002_s N_X_M1014_s
+ N_X_c_581_n N_X_c_582_n N_X_c_627_p N_X_c_578_n N_X_c_579_n N_X_c_615_n
+ N_X_c_583_n N_X_c_626_p N_X_c_619_n N_X_c_584_n X X X
+ PM_SKY130_FD_SC_LP__O22A_4%X
x_PM_SKY130_FD_SC_LP__O22A_4%A_608_367# N_A_608_367#_M1003_d
+ N_A_608_367#_M1018_d N_A_608_367#_c_634_n N_A_608_367#_c_635_n
+ N_A_608_367#_c_646_n N_A_608_367#_c_637_n
+ PM_SKY130_FD_SC_LP__O22A_4%A_608_367#
x_PM_SKY130_FD_SC_LP__O22A_4%A_982_367# N_A_982_367#_M1007_s
+ N_A_982_367#_M1017_s N_A_982_367#_c_649_n N_A_982_367#_c_650_n
+ N_A_982_367#_c_653_n N_A_982_367#_c_663_n N_A_982_367#_c_654_n
+ PM_SKY130_FD_SC_LP__O22A_4%A_982_367#
x_PM_SKY130_FD_SC_LP__O22A_4%VGND N_VGND_M1005_s N_VGND_M1011_s N_VGND_M1016_s
+ N_VGND_M1000_d N_VGND_M1020_d N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ N_VGND_c_668_n N_VGND_c_669_n N_VGND_c_670_n N_VGND_c_671_n N_VGND_c_672_n
+ N_VGND_c_673_n N_VGND_c_674_n VGND N_VGND_c_675_n N_VGND_c_676_n
+ N_VGND_c_677_n N_VGND_c_678_n N_VGND_c_679_n N_VGND_c_680_n
+ PM_SKY130_FD_SC_LP__O22A_4%VGND
x_PM_SKY130_FD_SC_LP__O22A_4%A_525_47# N_A_525_47#_M1010_s N_A_525_47#_M1006_s
+ N_A_525_47#_M1019_s N_A_525_47#_M1004_s N_A_525_47#_M1012_s
+ N_A_525_47#_c_768_n N_A_525_47#_c_805_n N_A_525_47#_c_787_n
+ N_A_525_47#_c_812_n N_A_525_47#_c_791_n N_A_525_47#_c_764_n
+ N_A_525_47#_c_765_n N_A_525_47#_c_770_n N_A_525_47#_c_782_n
+ N_A_525_47#_c_796_n PM_SKY130_FD_SC_LP__O22A_4%A_525_47#
cc_1 VNB N_A_86_23#_M1005_g 0.0266002f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.665
cc_2 VNB N_A_86_23#_M1011_g 0.0213855f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.665
cc_3 VNB N_A_86_23#_M1015_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.665
cc_4 VNB N_A_86_23#_M1016_g 0.0275234f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.665
cc_5 VNB N_A_86_23#_c_102_n 0.0179317f $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=1.405
cc_6 VNB N_A_86_23#_c_103_n 0.00470404f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=0.385
cc_7 VNB N_A_86_23#_c_104_n 0.00841275f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=0.4
cc_8 VNB N_A_86_23#_c_105_n 0.00120159f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=1.93
cc_9 VNB N_A_86_23#_c_106_n 0.00572131f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=1.49
cc_10 VNB N_A_86_23#_c_107_n 0.12057f $X=-0.19 $Y=-0.245 $X2=2.46 $Y2=1.49
cc_11 VNB N_B1_M1003_g 0.00727196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_M1023_g 0.00824325f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.325
cc_13 VNB N_B1_c_248_n 0.0156348f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.665
cc_14 VNB N_B1_c_249_n 0.0063608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_250_n 0.00335229f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.325
cc_16 VNB N_B1_c_251_n 0.032335f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.655
cc_17 VNB N_B1_c_252_n 0.0319142f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.665
cc_18 VNB N_B1_c_253_n 0.0200294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_254_n 0.0160938f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.465
cc_20 VNB N_B2_M1006_g 0.0226643f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=1.835
cc_21 VNB N_B2_M1021_g 0.0226358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B2_c_329_n 0.0326658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_M1007_g 0.00824313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_M1013_g 0.0080507f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.325
cc_25 VNB N_A1_c_374_n 0.0176407f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.665
cc_26 VNB N_A1_c_375_n 0.00338197f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.325
cc_27 VNB N_A1_c_376_n 0.0323294f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.655
cc_28 VNB A1 0.0313794f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.325
cc_29 VNB N_A1_c_378_n 0.0167172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_379_n 0.0356828f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.665
cc_31 VNB N_A1_c_380_n 0.0214439f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.655
cc_32 VNB N_A2_M1004_g 0.0232631f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=1.835
cc_33 VNB N_A2_M1020_g 0.0228415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB A2 0.00226109f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.325
cc_35 VNB N_A2_c_446_n 0.0316223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_490_n 0.283096f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.49
cc_37 VNB N_X_c_578_n 0.00663052f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.665
cc_38 VNB N_X_c_579_n 0.0129129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB X 0.020096f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.49
cc_40 VNB N_VGND_c_665_n 0.0113984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_666_n 0.0281531f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.665
cc_42 VNB N_VGND_c_667_n 4.82391e-19 $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=2.465
cc_43 VNB N_VGND_c_668_n 0.0070685f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.665
cc_44 VNB N_VGND_c_669_n 0.00496727f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.465
cc_45 VNB N_VGND_c_670_n 4.06069e-19 $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.665
cc_46 VNB N_VGND_c_671_n 0.014949f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.655
cc_47 VNB N_VGND_c_672_n 0.00461634f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.465
cc_48 VNB N_VGND_c_673_n 0.0136274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_674_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=2.46 $Y2=1.655
cc_50 VNB N_VGND_c_675_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_676_n 0.0639492f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=0.385
cc_52 VNB N_VGND_c_677_n 0.0185665f $X=-0.19 $Y=-0.245 $X2=3.775 $Y2=2.015
cc_53 VNB N_VGND_c_678_n 0.343342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_679_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_680_n 0.00632006f $X=-0.19 $Y=-0.245 $X2=5.48 $Y2=2.015
cc_56 VNB N_A_525_47#_c_764_n 0.0117193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_525_47#_c_765_n 0.0183124f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.665
cc_58 VPB N_A_86_23#_M1002_g 0.0232636f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.465
cc_59 VPB N_A_86_23#_M1009_g 0.0188632f $X=-0.19 $Y=1.655 $X2=1.6 $Y2=2.465
cc_60 VPB N_A_86_23#_M1014_g 0.0188559f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=2.465
cc_61 VPB N_A_86_23#_M1022_g 0.0199015f $X=-0.19 $Y=1.655 $X2=2.46 $Y2=2.465
cc_62 VPB N_A_86_23#_c_105_n 0.00177852f $X=-0.19 $Y=1.655 $X2=2.595 $Y2=1.93
cc_63 VPB N_A_86_23#_c_107_n 0.0242481f $X=-0.19 $Y=1.655 $X2=2.46 $Y2=1.49
cc_64 VPB N_B1_M1003_g 0.0213129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B1_M1023_g 0.02213f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.325
cc_66 VPB N_B2_M1008_g 0.018718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_B2_M1018_g 0.0187204f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.665
cc_68 VPB N_B2_c_332_n 0.00259388f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.465
cc_69 VPB N_B2_c_329_n 0.00488677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A1_M1007_g 0.02213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A1_M1013_g 0.0244984f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.325
cc_72 VPB A1 0.0172414f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=1.325
cc_73 VPB N_A2_M1001_g 0.0182421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A2_M1017_g 0.0186932f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.665
cc_75 VPB A2 0.0038254f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=1.325
cc_76 VPB N_A2_c_446_n 0.00474776f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_491_n 0.0414999f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.665
cc_78 VPB N_VPWR_c_492_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.465
cc_79 VPB N_VPWR_c_493_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.665
cc_80 VPB N_VPWR_c_494_n 0.00496093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_495_n 0.00557358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_496_n 0.0141676f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=2.465
cc_83 VPB N_VPWR_c_497_n 0.0476787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_498_n 0.0272827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_499_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.49
cc_86 VPB N_VPWR_c_500_n 0.0151004f $X=-0.19 $Y=1.655 $X2=2.465 $Y2=0.385
cc_87 VPB N_VPWR_c_501_n 0.0365476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_502_n 0.0346042f $X=-0.19 $Y=1.655 $X2=3.775 $Y2=2.015
cc_89 VPB N_VPWR_c_503_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.61 $Y2=2.095
cc_90 VPB N_VPWR_c_504_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.49
cc_91 VPB N_VPWR_c_505_n 0.00631788f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.49
cc_92 VPB N_VPWR_c_490_n 0.0778531f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=1.49
cc_93 VPB N_X_c_581_n 0.0162801f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.325
cc_94 VPB N_X_c_582_n 0.0258942f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.665
cc_95 VPB N_X_c_583_n 0.00512804f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.665
cc_96 VPB N_X_c_584_n 0.00147023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB X 0.00593595f $X=-0.19 $Y=1.655 $X2=0.94 $Y2=1.49
cc_98 N_A_86_23#_c_105_n N_B1_M1003_g 0.00723323f $X=2.595 $Y=1.93 $X2=0 $Y2=0
cc_99 N_A_86_23#_c_115_p N_B1_M1003_g 0.0166325f $X=3.445 $Y=2.015 $X2=0 $Y2=0
cc_100 N_A_86_23#_c_106_n N_B1_M1003_g 0.00131885f $X=2.595 $Y=1.49 $X2=0 $Y2=0
cc_101 N_A_86_23#_c_117_p N_B1_M1003_g 8.92984e-19 $X=3.61 $Y=2.095 $X2=0 $Y2=0
cc_102 N_A_86_23#_c_107_n N_B1_M1003_g 0.0303741f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_103 N_A_86_23#_c_119_p N_B1_M1023_g 0.0162758f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_104 N_A_86_23#_c_117_p N_B1_M1023_g 9.31581e-19 $X=3.61 $Y=2.095 $X2=0 $Y2=0
cc_105 N_A_86_23#_M1010_d N_B1_c_249_n 0.00268388f $X=3.04 $Y=0.235 $X2=0 $Y2=0
cc_106 N_A_86_23#_c_102_n N_B1_c_249_n 0.0121445f $X=2.38 $Y=1.405 $X2=0 $Y2=0
cc_107 N_A_86_23#_c_115_p N_B1_c_249_n 0.0146609f $X=3.445 $Y=2.015 $X2=0 $Y2=0
cc_108 N_A_86_23#_c_106_n N_B1_c_249_n 0.00982505f $X=2.595 $Y=1.49 $X2=0 $Y2=0
cc_109 N_A_86_23#_c_107_n N_B1_c_249_n 4.21722e-19 $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_110 N_A_86_23#_M1021_d N_B1_c_250_n 7.5535e-19 $X=3.9 $Y=0.235 $X2=0 $Y2=0
cc_111 N_A_86_23#_c_119_p N_B1_c_250_n 0.00996124f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_112 N_A_86_23#_c_119_p N_B1_c_251_n 6.72748e-19 $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_113 N_A_86_23#_c_102_n N_B1_c_252_n 0.00299255f $X=2.38 $Y=1.405 $X2=0 $Y2=0
cc_114 N_A_86_23#_c_115_p N_B1_c_252_n 0.00220882f $X=3.445 $Y=2.015 $X2=0 $Y2=0
cc_115 N_A_86_23#_c_106_n N_B1_c_252_n 9.24651e-19 $X=2.595 $Y=1.49 $X2=0 $Y2=0
cc_116 N_A_86_23#_c_107_n N_B1_c_252_n 0.0105625f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_117 N_A_86_23#_c_102_n N_B1_c_253_n 0.00741871f $X=2.38 $Y=1.405 $X2=0 $Y2=0
cc_118 N_A_86_23#_c_104_n N_B1_c_253_n 0.0129203f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_119 N_A_86_23#_c_104_n N_B1_c_254_n 0.00325378f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_120 N_A_86_23#_c_104_n N_B2_M1006_g 0.0100622f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_121 N_A_86_23#_c_115_p N_B2_M1008_g 0.0148906f $X=3.445 $Y=2.015 $X2=0 $Y2=0
cc_122 N_A_86_23#_c_117_p N_B2_M1008_g 0.0108226f $X=3.61 $Y=2.095 $X2=0 $Y2=0
cc_123 N_A_86_23#_c_104_n N_B2_M1021_g 0.0100622f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_124 N_A_86_23#_c_119_p N_B2_M1018_g 0.0110405f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_125 N_A_86_23#_c_117_p N_B2_M1018_g 0.0104106f $X=3.61 $Y=2.095 $X2=0 $Y2=0
cc_126 N_A_86_23#_c_119_p N_B2_c_332_n 0.00889924f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_127 N_A_86_23#_c_117_p N_B2_c_332_n 0.0223835f $X=3.61 $Y=2.095 $X2=0 $Y2=0
cc_128 N_A_86_23#_c_117_p N_B2_c_329_n 6.3648e-19 $X=3.61 $Y=2.095 $X2=0 $Y2=0
cc_129 N_A_86_23#_c_119_p N_A1_M1007_g 0.0162758f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_130 N_A_86_23#_c_146_p N_A1_M1007_g 9.31581e-19 $X=5.48 $Y=2.095 $X2=0 $Y2=0
cc_131 N_A_86_23#_c_119_p N_A1_c_375_n 0.00996124f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_132 N_A_86_23#_c_119_p N_A1_c_376_n 6.69142e-19 $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_133 N_A_86_23#_c_119_p N_A2_M1001_g 0.0111034f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_134 N_A_86_23#_c_146_p N_A2_M1001_g 0.0104718f $X=5.48 $Y=2.095 $X2=0 $Y2=0
cc_135 N_A_86_23#_c_146_p N_A2_M1017_g 0.0105296f $X=5.48 $Y=2.095 $X2=0 $Y2=0
cc_136 N_A_86_23#_c_119_p A2 0.00890349f $X=5.315 $Y=2.015 $X2=0 $Y2=0
cc_137 N_A_86_23#_c_146_p A2 0.0230948f $X=5.48 $Y=2.095 $X2=0 $Y2=0
cc_138 N_A_86_23#_c_146_p N_A2_c_446_n 6.37898e-19 $X=5.48 $Y=2.095 $X2=0 $Y2=0
cc_139 N_A_86_23#_c_105_n N_VPWR_M1022_d 0.00112177f $X=2.595 $Y=1.93 $X2=0
+ $Y2=0
cc_140 N_A_86_23#_c_115_p N_VPWR_M1022_d 0.00614282f $X=3.445 $Y=2.015 $X2=0
+ $Y2=0
cc_141 N_A_86_23#_c_157_p N_VPWR_M1022_d 9.55196e-19 $X=2.68 $Y=2.015 $X2=0
+ $Y2=0
cc_142 N_A_86_23#_c_119_p N_VPWR_M1023_s 0.0135034f $X=5.315 $Y=2.015 $X2=0
+ $Y2=0
cc_143 N_A_86_23#_M1002_g N_VPWR_c_491_n 0.0152824f $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_86_23#_M1009_g N_VPWR_c_491_n 7.27171e-19 $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_86_23#_M1002_g N_VPWR_c_492_n 0.00486043f $X=1.17 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_86_23#_M1009_g N_VPWR_c_492_n 0.00486043f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_86_23#_M1002_g N_VPWR_c_493_n 7.24342e-19 $X=1.17 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_86_23#_M1009_g N_VPWR_c_493_n 0.0141279f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_86_23#_M1014_g N_VPWR_c_493_n 0.0142085f $X=2.03 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_86_23#_M1022_g N_VPWR_c_493_n 7.38561e-19 $X=2.46 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_86_23#_M1022_g N_VPWR_c_494_n 0.00261698f $X=2.46 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_86_23#_c_115_p N_VPWR_c_494_n 0.0124114f $X=3.445 $Y=2.015 $X2=0
+ $Y2=0
cc_153 N_A_86_23#_c_157_p N_VPWR_c_494_n 0.00774152f $X=2.68 $Y=2.015 $X2=0
+ $Y2=0
cc_154 N_A_86_23#_c_119_p N_VPWR_c_495_n 0.0257093f $X=5.315 $Y=2.015 $X2=0
+ $Y2=0
cc_155 N_A_86_23#_M1014_g N_VPWR_c_500_n 0.00486043f $X=2.03 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_86_23#_M1022_g N_VPWR_c_500_n 0.00585385f $X=2.46 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_86_23#_M1008_s N_VPWR_c_490_n 0.00225186f $X=3.47 $Y=1.835 $X2=0
+ $Y2=0
cc_158 N_A_86_23#_M1001_d N_VPWR_c_490_n 0.00225186f $X=5.34 $Y=1.835 $X2=0
+ $Y2=0
cc_159 N_A_86_23#_M1002_g N_VPWR_c_490_n 0.00824727f $X=1.17 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_86_23#_M1009_g N_VPWR_c_490_n 0.00824727f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A_86_23#_M1014_g N_VPWR_c_490_n 0.00824727f $X=2.03 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_86_23#_M1022_g N_VPWR_c_490_n 0.010718f $X=2.46 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_86_23#_M1002_g N_X_c_581_n 0.0153141f $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A_86_23#_c_180_p N_X_c_581_n 0.0346829f $X=2.295 $Y=1.49 $X2=0 $Y2=0
cc_165 N_A_86_23#_c_107_n N_X_c_581_n 0.0176339f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_166 N_A_86_23#_M1011_g N_X_c_578_n 0.0139493f $X=0.935 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A_86_23#_M1015_g N_X_c_578_n 0.013726f $X=1.365 $Y=0.665 $X2=0 $Y2=0
cc_168 N_A_86_23#_M1016_g N_X_c_578_n 0.00219965f $X=1.795 $Y=0.665 $X2=0 $Y2=0
cc_169 N_A_86_23#_c_180_p N_X_c_578_n 0.0177796f $X=2.295 $Y=1.49 $X2=0 $Y2=0
cc_170 N_A_86_23#_c_102_n N_X_c_578_n 0.00426737f $X=2.38 $Y=1.405 $X2=0 $Y2=0
cc_171 N_A_86_23#_c_107_n N_X_c_578_n 0.00585496f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_172 N_A_86_23#_M1005_g N_X_c_579_n 0.0152898f $X=0.505 $Y=0.665 $X2=0 $Y2=0
cc_173 N_A_86_23#_c_180_p N_X_c_579_n 0.0474479f $X=2.295 $Y=1.49 $X2=0 $Y2=0
cc_174 N_A_86_23#_c_107_n N_X_c_579_n 0.0028595f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_175 N_A_86_23#_M1009_g N_X_c_583_n 0.0132368f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_86_23#_M1014_g N_X_c_583_n 0.0130747f $X=2.03 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A_86_23#_M1022_g N_X_c_583_n 6.55961e-19 $X=2.46 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_86_23#_c_180_p N_X_c_583_n 0.0593284f $X=2.295 $Y=1.49 $X2=0 $Y2=0
cc_179 N_A_86_23#_c_105_n N_X_c_583_n 0.00947164f $X=2.595 $Y=1.93 $X2=0 $Y2=0
cc_180 N_A_86_23#_c_107_n N_X_c_583_n 0.00542936f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_181 N_A_86_23#_c_180_p N_X_c_584_n 0.014687f $X=2.295 $Y=1.49 $X2=0 $Y2=0
cc_182 N_A_86_23#_c_107_n N_X_c_584_n 0.00298081f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_183 N_A_86_23#_M1005_g X 0.00452206f $X=0.505 $Y=0.665 $X2=0 $Y2=0
cc_184 N_A_86_23#_M1011_g X 5.295e-19 $X=0.935 $Y=0.665 $X2=0 $Y2=0
cc_185 N_A_86_23#_M1002_g X 0.00244719f $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_86_23#_c_180_p X 0.00941438f $X=2.295 $Y=1.49 $X2=0 $Y2=0
cc_187 N_A_86_23#_c_107_n X 0.0216244f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_188 N_A_86_23#_c_115_p N_A_608_367#_M1003_d 0.00440504f $X=3.445 $Y=2.015
+ $X2=-0.19 $Y2=-0.245
cc_189 N_A_86_23#_c_119_p N_A_608_367#_M1018_d 0.0078026f $X=5.315 $Y=2.015
+ $X2=0 $Y2=0
cc_190 N_A_86_23#_c_115_p N_A_608_367#_c_634_n 0.0135055f $X=3.445 $Y=2.015
+ $X2=0 $Y2=0
cc_191 N_A_86_23#_M1008_s N_A_608_367#_c_635_n 0.00332344f $X=3.47 $Y=1.835
+ $X2=0 $Y2=0
cc_192 N_A_86_23#_c_117_p N_A_608_367#_c_635_n 0.0159805f $X=3.61 $Y=2.095 $X2=0
+ $Y2=0
cc_193 N_A_86_23#_c_119_p N_A_608_367#_c_637_n 0.0152916f $X=5.315 $Y=2.015
+ $X2=0 $Y2=0
cc_194 N_A_86_23#_c_119_p N_A_982_367#_M1007_s 0.0078026f $X=5.315 $Y=2.015
+ $X2=-0.19 $Y2=-0.245
cc_195 N_A_86_23#_c_119_p N_A_982_367#_c_649_n 0.0152916f $X=5.315 $Y=2.015
+ $X2=0 $Y2=0
cc_196 N_A_86_23#_M1001_d N_A_982_367#_c_650_n 0.00332344f $X=5.34 $Y=1.835
+ $X2=0 $Y2=0
cc_197 N_A_86_23#_c_146_p N_A_982_367#_c_650_n 0.0159805f $X=5.48 $Y=2.095 $X2=0
+ $Y2=0
cc_198 N_A_86_23#_M1005_g N_VGND_c_666_n 0.0116205f $X=0.505 $Y=0.665 $X2=0
+ $Y2=0
cc_199 N_A_86_23#_M1011_g N_VGND_c_666_n 6.10117e-19 $X=0.935 $Y=0.665 $X2=0
+ $Y2=0
cc_200 N_A_86_23#_M1005_g N_VGND_c_667_n 6.10117e-19 $X=0.505 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_86_23#_M1011_g N_VGND_c_667_n 0.0107978f $X=0.935 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_86_23#_M1015_g N_VGND_c_667_n 0.0108835f $X=1.365 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_86_23#_M1016_g N_VGND_c_667_n 6.25217e-19 $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_204 N_A_86_23#_M1016_g N_VGND_c_668_n 0.00696134f $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_205 N_A_86_23#_c_180_p N_VGND_c_668_n 0.0125999f $X=2.295 $Y=1.49 $X2=0 $Y2=0
cc_206 N_A_86_23#_c_102_n N_VGND_c_668_n 0.0447667f $X=2.38 $Y=1.405 $X2=0 $Y2=0
cc_207 N_A_86_23#_c_103_n N_VGND_c_668_n 0.0221159f $X=2.465 $Y=0.385 $X2=0
+ $Y2=0
cc_208 N_A_86_23#_c_107_n N_VGND_c_668_n 0.00655957f $X=2.46 $Y=1.49 $X2=0 $Y2=0
cc_209 N_A_86_23#_M1015_g N_VGND_c_671_n 0.00477554f $X=1.365 $Y=0.665 $X2=0
+ $Y2=0
cc_210 N_A_86_23#_M1016_g N_VGND_c_671_n 0.00575161f $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_86_23#_M1005_g N_VGND_c_675_n 0.00477554f $X=0.505 $Y=0.665 $X2=0
+ $Y2=0
cc_212 N_A_86_23#_M1011_g N_VGND_c_675_n 0.00477554f $X=0.935 $Y=0.665 $X2=0
+ $Y2=0
cc_213 N_A_86_23#_c_103_n N_VGND_c_676_n 0.0121867f $X=2.465 $Y=0.385 $X2=0
+ $Y2=0
cc_214 N_A_86_23#_c_104_n N_VGND_c_676_n 0.100659f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_215 N_A_86_23#_M1010_d N_VGND_c_678_n 0.00223577f $X=3.04 $Y=0.235 $X2=0
+ $Y2=0
cc_216 N_A_86_23#_M1021_d N_VGND_c_678_n 0.00223577f $X=3.9 $Y=0.235 $X2=0 $Y2=0
cc_217 N_A_86_23#_M1005_g N_VGND_c_678_n 0.00825815f $X=0.505 $Y=0.665 $X2=0
+ $Y2=0
cc_218 N_A_86_23#_M1011_g N_VGND_c_678_n 0.00825815f $X=0.935 $Y=0.665 $X2=0
+ $Y2=0
cc_219 N_A_86_23#_M1015_g N_VGND_c_678_n 0.00825815f $X=1.365 $Y=0.665 $X2=0
+ $Y2=0
cc_220 N_A_86_23#_M1016_g N_VGND_c_678_n 0.0118487f $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_221 N_A_86_23#_c_103_n N_VGND_c_678_n 0.00660921f $X=2.465 $Y=0.385 $X2=0
+ $Y2=0
cc_222 N_A_86_23#_c_104_n N_VGND_c_678_n 0.0635746f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_223 N_A_86_23#_c_104_n N_A_525_47#_M1010_s 0.00569291f $X=4.04 $Y=0.4
+ $X2=-0.19 $Y2=-0.245
cc_224 N_A_86_23#_c_104_n N_A_525_47#_M1006_s 0.0033716f $X=4.04 $Y=0.4 $X2=0
+ $Y2=0
cc_225 N_A_86_23#_M1010_d N_A_525_47#_c_768_n 0.00348247f $X=3.04 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_A_86_23#_M1021_d N_A_525_47#_c_768_n 0.00347723f $X=3.9 $Y=0.235 $X2=0
+ $Y2=0
cc_227 N_A_86_23#_c_102_n N_A_525_47#_c_770_n 0.0263952f $X=2.38 $Y=1.405 $X2=0
+ $Y2=0
cc_228 N_A_86_23#_c_104_n N_A_525_47#_c_770_n 0.0835599f $X=4.04 $Y=0.4 $X2=0
+ $Y2=0
cc_229 N_A_86_23#_c_106_n N_A_525_47#_c_770_n 0.00193438f $X=2.595 $Y=1.49 $X2=0
+ $Y2=0
cc_230 N_B1_c_248_n N_B2_M1006_g 0.0144197f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B1_c_249_n N_B2_M1006_g 0.00578897f $X=3.285 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B1_c_252_n N_B2_M1006_g 0.020614f $X=2.945 $Y=1.36 $X2=0 $Y2=0
cc_233 N_B1_c_253_n N_B2_M1006_g 0.0345333f $X=2.945 $Y=1.195 $X2=0 $Y2=0
cc_234 N_B1_c_248_n N_B2_M1021_g 0.00995077f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B1_c_250_n N_B2_M1021_g 0.00171593f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B1_c_251_n N_B2_M1021_g 0.0215587f $X=4.275 $Y=1.35 $X2=0 $Y2=0
cc_237 N_B1_c_254_n N_B2_M1021_g 0.0341982f $X=4.275 $Y=1.185 $X2=0 $Y2=0
cc_238 N_B1_M1003_g N_B2_c_332_n 0.00111536f $X=2.965 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1023_g N_B2_c_332_n 0.00152269f $X=4.255 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_c_248_n N_B2_c_332_n 0.0329645f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_241 N_B1_c_249_n N_B2_c_332_n 0.00911937f $X=3.285 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B1_c_250_n N_B2_c_332_n 0.00648564f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B1_c_251_n N_B2_c_332_n 3.47814e-19 $X=4.275 $Y=1.35 $X2=0 $Y2=0
cc_244 N_B1_M1003_g N_B2_c_329_n 0.0423567f $X=2.965 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_M1023_g N_B2_c_329_n 0.044384f $X=4.255 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B1_c_248_n N_B2_c_329_n 0.00243405f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_247 N_B1_M1023_g N_A1_M1007_g 0.0435212f $X=4.255 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B1_c_250_n N_A1_c_375_n 0.0288098f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_249 N_B1_c_251_n N_A1_c_375_n 0.00114936f $X=4.275 $Y=1.35 $X2=0 $Y2=0
cc_250 N_B1_c_254_n N_A1_c_375_n 3.35101e-19 $X=4.275 $Y=1.185 $X2=0 $Y2=0
cc_251 N_B1_c_250_n N_A1_c_376_n 0.00114936f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B1_c_251_n N_A1_c_376_n 0.0201104f $X=4.275 $Y=1.35 $X2=0 $Y2=0
cc_253 N_B1_c_250_n N_A1_c_378_n 3.90691e-19 $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B1_c_254_n N_A1_c_378_n 0.0223037f $X=4.275 $Y=1.185 $X2=0 $Y2=0
cc_255 N_B1_M1003_g N_VPWR_c_494_n 0.00413277f $X=2.965 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B1_M1023_g N_VPWR_c_495_n 0.0081983f $X=4.255 $Y=2.465 $X2=0 $Y2=0
cc_257 N_B1_M1003_g N_VPWR_c_501_n 0.00585385f $X=2.965 $Y=2.465 $X2=0 $Y2=0
cc_258 N_B1_M1023_g N_VPWR_c_501_n 0.00547432f $X=4.255 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B1_M1003_g N_VPWR_c_490_n 0.010757f $X=2.965 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B1_M1023_g N_VPWR_c_490_n 0.0102457f $X=4.255 $Y=2.465 $X2=0 $Y2=0
cc_261 N_B1_M1023_g N_A_608_367#_c_635_n 0.0019889f $X=4.255 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_B1_M1023_g N_A_608_367#_c_637_n 0.00775016f $X=4.255 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_B1_c_253_n N_VGND_c_676_n 0.00357877f $X=2.945 $Y=1.195 $X2=0 $Y2=0
cc_264 N_B1_c_254_n N_VGND_c_676_n 0.00419907f $X=4.275 $Y=1.185 $X2=0 $Y2=0
cc_265 N_B1_c_253_n N_VGND_c_678_n 0.0067762f $X=2.945 $Y=1.195 $X2=0 $Y2=0
cc_266 N_B1_c_254_n N_VGND_c_678_n 0.00620263f $X=4.275 $Y=1.185 $X2=0 $Y2=0
cc_267 N_B1_c_250_n N_A_525_47#_M1019_s 0.00119179f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_268 N_B1_c_248_n N_A_525_47#_c_768_n 0.052445f $X=4.11 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B1_c_249_n N_A_525_47#_c_768_n 0.0245115f $X=3.285 $Y=1.16 $X2=0 $Y2=0
cc_270 N_B1_c_250_n N_A_525_47#_c_768_n 0.0169002f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B1_c_251_n N_A_525_47#_c_768_n 2.67964e-19 $X=4.275 $Y=1.35 $X2=0 $Y2=0
cc_272 N_B1_c_252_n N_A_525_47#_c_768_n 2.67022e-19 $X=2.945 $Y=1.36 $X2=0 $Y2=0
cc_273 N_B1_c_253_n N_A_525_47#_c_768_n 0.0103716f $X=2.945 $Y=1.195 $X2=0 $Y2=0
cc_274 N_B1_c_254_n N_A_525_47#_c_768_n 0.0140999f $X=4.275 $Y=1.185 $X2=0 $Y2=0
cc_275 N_B1_c_252_n N_A_525_47#_c_770_n 0.00265979f $X=2.945 $Y=1.36 $X2=0 $Y2=0
cc_276 N_B1_c_250_n N_A_525_47#_c_782_n 0.0046107f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_277 N_B1_c_251_n N_A_525_47#_c_782_n 3.16955e-19 $X=4.275 $Y=1.35 $X2=0 $Y2=0
cc_278 N_B2_M1008_g N_VPWR_c_501_n 0.00357877f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_279 N_B2_M1018_g N_VPWR_c_501_n 0.00357877f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_280 N_B2_M1008_g N_VPWR_c_490_n 0.00537654f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_281 N_B2_M1018_g N_VPWR_c_490_n 0.00537654f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_282 N_B2_M1008_g N_A_608_367#_c_635_n 0.0115031f $X=3.395 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_B2_M1018_g N_A_608_367#_c_635_n 0.0114565f $X=3.825 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_B2_M1006_g N_VGND_c_676_n 0.00357877f $X=3.395 $Y=0.655 $X2=0 $Y2=0
cc_285 N_B2_M1021_g N_VGND_c_676_n 0.00357877f $X=3.825 $Y=0.655 $X2=0 $Y2=0
cc_286 N_B2_M1006_g N_VGND_c_678_n 0.00537654f $X=3.395 $Y=0.655 $X2=0 $Y2=0
cc_287 N_B2_M1021_g N_VGND_c_678_n 0.00537654f $X=3.825 $Y=0.655 $X2=0 $Y2=0
cc_288 N_B2_M1006_g N_A_525_47#_c_768_n 0.00970969f $X=3.395 $Y=0.655 $X2=0
+ $Y2=0
cc_289 N_B2_M1021_g N_A_525_47#_c_768_n 0.00969584f $X=3.825 $Y=0.655 $X2=0
+ $Y2=0
cc_290 N_A1_c_374_n N_A2_M1004_g 0.0101984f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A1_c_375_n N_A2_M1004_g 0.00143125f $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A1_c_376_n N_A2_M1004_g 0.0215822f $X=4.815 $Y=1.35 $X2=0 $Y2=0
cc_293 N_A1_c_378_n N_A2_M1004_g 0.0251033f $X=4.815 $Y=1.185 $X2=0 $Y2=0
cc_294 N_A1_c_374_n N_A2_M1020_g 0.0131727f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_295 A1 N_A2_M1020_g 0.00890876f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_296 N_A1_c_380_n N_A2_M1020_g 0.0237068f $X=6.215 $Y=1.185 $X2=0 $Y2=0
cc_297 N_A1_M1013_g N_A2_M1017_g 0.0237068f $X=6.125 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A1_M1007_g A2 0.0015176f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A1_c_374_n A2 0.0345242f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A1_c_375_n A2 0.00584007f $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A1_c_376_n A2 3.09875e-19 $X=4.815 $Y=1.35 $X2=0 $Y2=0
cc_302 A1 A2 0.0289592f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_303 N_A1_c_379_n A2 2.67103e-19 $X=6.215 $Y=1.35 $X2=0 $Y2=0
cc_304 N_A1_M1007_g N_A2_c_446_n 0.0428136f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A1_c_374_n N_A2_c_446_n 0.00244902f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A1_c_379_n N_A2_c_446_n 0.0237068f $X=6.215 $Y=1.35 $X2=0 $Y2=0
cc_307 N_A1_M1007_g N_VPWR_c_495_n 0.0081983f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A1_M1013_g N_VPWR_c_497_n 0.0209615f $X=6.125 $Y=2.465 $X2=0 $Y2=0
cc_309 A1 N_VPWR_c_497_n 0.0270936f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_310 N_A1_c_379_n N_VPWR_c_497_n 7.02047e-19 $X=6.215 $Y=1.35 $X2=0 $Y2=0
cc_311 N_A1_M1007_g N_VPWR_c_502_n 0.00547432f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A1_M1013_g N_VPWR_c_502_n 0.00486043f $X=6.125 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A1_M1007_g N_VPWR_c_490_n 0.0102457f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A1_M1013_g N_VPWR_c_490_n 0.0082726f $X=6.125 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A1_M1007_g N_A_982_367#_c_649_n 0.00775016f $X=4.835 $Y=2.465 $X2=0
+ $Y2=0
cc_316 N_A1_M1007_g N_A_982_367#_c_653_n 0.0019889f $X=4.835 $Y=2.465 $X2=0
+ $Y2=0
cc_317 A1 N_A_982_367#_c_654_n 0.013685f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_318 N_A1_c_375_n N_VGND_M1000_d 0.00152165f $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_319 A1 N_VGND_M1020_d 0.00222017f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_320 N_A1_c_378_n N_VGND_c_669_n 0.00336962f $X=4.815 $Y=1.185 $X2=0 $Y2=0
cc_321 N_A1_c_380_n N_VGND_c_670_n 0.00909689f $X=6.215 $Y=1.185 $X2=0 $Y2=0
cc_322 N_A1_c_378_n N_VGND_c_676_n 0.00439206f $X=4.815 $Y=1.185 $X2=0 $Y2=0
cc_323 N_A1_c_380_n N_VGND_c_677_n 0.00365202f $X=6.215 $Y=1.185 $X2=0 $Y2=0
cc_324 N_A1_c_378_n N_VGND_c_678_n 0.00632833f $X=4.815 $Y=1.185 $X2=0 $Y2=0
cc_325 N_A1_c_380_n N_VGND_c_678_n 0.00535042f $X=6.215 $Y=1.185 $X2=0 $Y2=0
cc_326 N_A1_c_375_n N_A_525_47#_M1019_s 4.26293e-19 $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A1_c_374_n N_A_525_47#_c_787_n 0.0237845f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A1_c_375_n N_A_525_47#_c_787_n 0.0204579f $X=4.815 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A1_c_376_n N_A_525_47#_c_787_n 6.34307e-19 $X=4.815 $Y=1.35 $X2=0 $Y2=0
cc_330 N_A1_c_378_n N_A_525_47#_c_787_n 0.0105408f $X=4.815 $Y=1.185 $X2=0 $Y2=0
cc_331 N_A1_c_374_n N_A_525_47#_c_791_n 0.0156371f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_332 A1 N_A_525_47#_c_791_n 0.0225765f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_333 N_A1_c_380_n N_A_525_47#_c_791_n 0.0104566f $X=6.215 $Y=1.185 $X2=0 $Y2=0
cc_334 A1 N_A_525_47#_c_764_n 0.0233876f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_335 N_A1_c_379_n N_A_525_47#_c_764_n 0.00112981f $X=6.215 $Y=1.35 $X2=0 $Y2=0
cc_336 N_A1_c_374_n N_A_525_47#_c_796_n 0.0160965f $X=5.85 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A2_M1017_g N_VPWR_c_497_n 0.00109252f $X=5.695 $Y=2.465 $X2=0 $Y2=0
cc_338 N_A2_M1001_g N_VPWR_c_502_n 0.00357877f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A2_M1017_g N_VPWR_c_502_n 0.00357877f $X=5.695 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A2_M1001_g N_VPWR_c_490_n 0.00537654f $X=5.265 $Y=2.465 $X2=0 $Y2=0
cc_341 N_A2_M1017_g N_VPWR_c_490_n 0.00537654f $X=5.695 $Y=2.465 $X2=0 $Y2=0
cc_342 N_A2_M1001_g N_A_982_367#_c_650_n 0.0114565f $X=5.265 $Y=2.465 $X2=0
+ $Y2=0
cc_343 N_A2_M1017_g N_A_982_367#_c_650_n 0.0115031f $X=5.695 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A2_M1004_g N_VGND_c_669_n 0.00176318f $X=5.265 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A2_M1004_g N_VGND_c_670_n 5.53848e-19 $X=5.265 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A2_M1020_g N_VGND_c_670_n 0.00763343f $X=5.695 $Y=0.655 $X2=0 $Y2=0
cc_347 N_A2_M1004_g N_VGND_c_673_n 0.00439206f $X=5.265 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A2_M1020_g N_VGND_c_673_n 0.00365202f $X=5.695 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A2_M1004_g N_VGND_c_678_n 0.00614948f $X=5.265 $Y=0.655 $X2=0 $Y2=0
cc_350 N_A2_M1020_g N_VGND_c_678_n 0.00432244f $X=5.695 $Y=0.655 $X2=0 $Y2=0
cc_351 N_A2_M1004_g N_A_525_47#_c_787_n 0.0105469f $X=5.265 $Y=0.655 $X2=0 $Y2=0
cc_352 N_A2_M1020_g N_A_525_47#_c_791_n 0.0098539f $X=5.695 $Y=0.655 $X2=0 $Y2=0
cc_353 N_VPWR_c_490_n N_X_M1002_s 0.00536646f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPWR_c_490_n N_X_M1014_s 0.00536646f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_355 N_VPWR_M1002_d N_X_c_581_n 0.00262981f $X=0.83 $Y=1.835 $X2=0 $Y2=0
cc_356 N_VPWR_c_491_n N_X_c_581_n 0.0220025f $X=0.955 $Y=2.18 $X2=0 $Y2=0
cc_357 N_VPWR_c_492_n N_X_c_615_n 0.0124525f $X=1.65 $Y=3.33 $X2=0 $Y2=0
cc_358 N_VPWR_c_490_n N_X_c_615_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_359 N_VPWR_M1009_d N_X_c_583_n 0.00180746f $X=1.675 $Y=1.835 $X2=0 $Y2=0
cc_360 N_VPWR_c_493_n N_X_c_583_n 0.0163515f $X=1.815 $Y=2.19 $X2=0 $Y2=0
cc_361 N_VPWR_c_500_n N_X_c_619_n 0.0124525f $X=2.545 $Y=3.33 $X2=0 $Y2=0
cc_362 N_VPWR_c_490_n N_X_c_619_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_363 N_VPWR_c_490_n N_A_608_367#_M1003_d 0.00220345f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_364 N_VPWR_c_490_n N_A_608_367#_M1018_d 0.00223562f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_501_n N_A_608_367#_c_635_n 0.0519089f $X=4.38 $Y=3.33 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_490_n N_A_608_367#_c_635_n 0.0335966f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_501_n N_A_608_367#_c_646_n 0.0139427f $X=4.38 $Y=3.33 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_490_n N_A_608_367#_c_646_n 0.00894187f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_490_n N_A_982_367#_M1007_s 0.00223562f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_370 N_VPWR_c_490_n N_A_982_367#_M1017_s 0.00376627f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_502_n N_A_982_367#_c_650_n 0.0361172f $X=6.175 $Y=3.33 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_490_n N_A_982_367#_c_650_n 0.023676f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_373 N_VPWR_c_502_n N_A_982_367#_c_653_n 0.0157917f $X=6.175 $Y=3.33 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_490_n N_A_982_367#_c_653_n 0.00992063f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_502_n N_A_982_367#_c_663_n 0.0125234f $X=6.175 $Y=3.33 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_490_n N_A_982_367#_c_663_n 0.00738676f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_377 N_X_c_579_n N_VGND_M1005_s 0.00234752f $X=0.815 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_378 N_X_c_578_n N_VGND_M1011_s 0.00176461f $X=1.485 $Y=1.14 $X2=0 $Y2=0
cc_379 N_X_c_579_n N_VGND_c_666_n 0.0220026f $X=0.815 $Y=1.14 $X2=0 $Y2=0
cc_380 N_X_c_578_n N_VGND_c_667_n 0.0170777f $X=1.485 $Y=1.14 $X2=0 $Y2=0
cc_381 N_X_c_578_n N_VGND_c_668_n 0.00164217f $X=1.485 $Y=1.14 $X2=0 $Y2=0
cc_382 N_X_c_626_p N_VGND_c_671_n 0.0138717f $X=1.58 $Y=0.42 $X2=0 $Y2=0
cc_383 N_X_c_627_p N_VGND_c_675_n 0.0124525f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_384 N_X_M1005_d N_VGND_c_678_n 0.00536646f $X=0.58 $Y=0.245 $X2=0 $Y2=0
cc_385 N_X_M1015_d N_VGND_c_678_n 0.00397496f $X=1.44 $Y=0.245 $X2=0 $Y2=0
cc_386 N_X_c_627_p N_VGND_c_678_n 0.00730901f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_387 N_X_c_626_p N_VGND_c_678_n 0.00886411f $X=1.58 $Y=0.42 $X2=0 $Y2=0
cc_388 N_VGND_c_678_n N_A_525_47#_M1010_s 0.0021598f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_389 N_VGND_c_678_n N_A_525_47#_M1006_s 0.00225186f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_678_n N_A_525_47#_M1019_s 0.00317914f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_c_678_n N_A_525_47#_M1004_s 0.00240997f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_678_n N_A_525_47#_M1012_s 0.00236587f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_676_n N_A_525_47#_c_768_n 0.00232518f $X=4.845 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_c_676_n N_A_525_47#_c_805_n 0.0187299f $X=4.845 $Y=0 $X2=0 $Y2=0
cc_395 N_VGND_c_678_n N_A_525_47#_c_805_n 0.0111782f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_M1000_d N_A_525_47#_c_787_n 0.00479363f $X=4.84 $Y=0.235 $X2=0
+ $Y2=0
cc_397 N_VGND_c_669_n N_A_525_47#_c_787_n 0.0185079f $X=5.01 $Y=0.44 $X2=0 $Y2=0
cc_398 N_VGND_c_673_n N_A_525_47#_c_787_n 0.00210007f $X=5.745 $Y=0 $X2=0 $Y2=0
cc_399 N_VGND_c_676_n N_A_525_47#_c_787_n 0.00210007f $X=4.845 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_678_n N_A_525_47#_c_787_n 0.00853765f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_673_n N_A_525_47#_c_812_n 0.0138332f $X=5.745 $Y=0 $X2=0 $Y2=0
cc_402 N_VGND_c_678_n N_A_525_47#_c_812_n 0.00885359f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_403 N_VGND_M1020_d N_A_525_47#_c_791_n 0.00348805f $X=5.77 $Y=0.235 $X2=0
+ $Y2=0
cc_404 N_VGND_c_670_n N_A_525_47#_c_791_n 0.016459f $X=5.91 $Y=0.44 $X2=0 $Y2=0
cc_405 N_VGND_c_673_n N_A_525_47#_c_791_n 0.00196209f $X=5.745 $Y=0 $X2=0 $Y2=0
cc_406 N_VGND_c_677_n N_A_525_47#_c_791_n 0.00181088f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_407 N_VGND_c_678_n N_A_525_47#_c_791_n 0.00838734f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_678_n N_A_525_47#_c_764_n 5.40712e-19 $X=6.48 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_677_n N_A_525_47#_c_765_n 0.0178111f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_678_n N_A_525_47#_c_765_n 0.0100304f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_678_n N_A_525_47#_c_770_n 0.00719861f $X=6.48 $Y=0 $X2=0 $Y2=0
