* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o31a_lp A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_37_57# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VGND a_37_57# a_516_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_37_57# B1 a_140_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_360_410# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VGND A2 a_140_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR B1 a_37_57# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_140_57# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_140_57# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_256_410# A2 a_360_410# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_516_57# a_37_57# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_37_57# A3 a_256_410# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
