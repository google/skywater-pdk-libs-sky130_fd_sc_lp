# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a221oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.830000 1.200000 8.075000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.410000 1.345000 6.660000 1.615000 ;
        RECT 6.410000 1.615000 8.485000 1.785000 ;
        RECT 8.245000 1.210000 9.995000 1.435000 ;
        RECT 8.245000 1.435000 8.485000 1.615000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.355000 5.680000 1.760000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805000 1.425000 3.815000 1.625000 ;
        RECT 3.645000 1.625000 3.815000 1.930000 ;
        RECT 3.645000 1.930000 6.085000 2.100000 ;
        RECT 5.850000 1.345000 6.200000 1.675000 ;
        RECT 5.850000 1.675000 6.085000 1.930000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 2.265000 1.435000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.116800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815000 1.605000 2.635000 1.775000 ;
        RECT 0.815000 1.775000 1.145000 2.735000 ;
        RECT 1.055000 0.255000 1.245000 0.870000 ;
        RECT 1.055000 0.870000 2.605000 1.015000 ;
        RECT 1.055000 1.015000 8.255000 1.030000 ;
        RECT 1.055000 1.030000 5.605000 1.040000 ;
        RECT 1.675000 1.775000 2.005000 2.735000 ;
        RECT 1.915000 0.255000 2.105000 0.870000 ;
        RECT 2.435000 1.040000 5.605000 1.185000 ;
        RECT 2.435000 1.185000 3.815000 1.255000 ;
        RECT 2.435000 1.255000 2.635000 1.605000 ;
        RECT 3.985000 0.755000 5.965000 0.860000 ;
        RECT 3.985000 0.860000 8.255000 1.015000 ;
        RECT 7.075000 0.700000 8.255000 0.860000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 10.080000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 10.270000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.385000  1.815000  0.645000 2.905000 ;
      RECT 0.385000  2.905000  2.435000 3.075000 ;
      RECT 0.555000  0.085000  0.885000 1.040000 ;
      RECT 1.315000  1.945000  1.505000 2.905000 ;
      RECT 1.415000  0.085000  1.745000 0.700000 ;
      RECT 2.175000  1.945000  3.325000 2.115000 ;
      RECT 2.175000  2.115000  2.435000 2.905000 ;
      RECT 2.275000  0.085000  2.605000 0.700000 ;
      RECT 2.625000  2.285000  2.955000 2.770000 ;
      RECT 2.625000  2.770000  6.455000 3.075000 ;
      RECT 2.775000  0.505000  2.965000 0.675000 ;
      RECT 2.775000  0.675000  3.815000 0.845000 ;
      RECT 3.055000  1.795000  3.325000 1.945000 ;
      RECT 3.125000  2.115000  3.325000 2.270000 ;
      RECT 3.125000  2.270000  5.965000 2.600000 ;
      RECT 3.135000  0.085000  3.465000 0.505000 ;
      RECT 3.635000  0.255000  5.955000 0.585000 ;
      RECT 3.635000  0.585000  3.815000 0.675000 ;
      RECT 6.135000  0.085000  6.465000 0.690000 ;
      RECT 6.135000  2.270000  6.455000 2.770000 ;
      RECT 6.255000  1.955000  9.055000 2.125000 ;
      RECT 6.255000  2.125000  6.455000 2.270000 ;
      RECT 6.625000  2.295000  6.955000 3.245000 ;
      RECT 6.645000  0.255000  8.625000 0.530000 ;
      RECT 7.135000  2.125000  7.335000 3.075000 ;
      RECT 7.505000  2.295000  7.835000 3.245000 ;
      RECT 8.005000  2.125000  8.195000 3.075000 ;
      RECT 8.365000  2.295000  8.695000 3.245000 ;
      RECT 8.425000  0.530000  8.625000 0.870000 ;
      RECT 8.425000  0.870000  9.485000 1.040000 ;
      RECT 8.795000  0.085000  9.125000 0.700000 ;
      RECT 8.795000  1.605000  9.985000 1.775000 ;
      RECT 8.795000  1.775000  9.055000 1.955000 ;
      RECT 8.865000  2.125000  9.055000 3.075000 ;
      RECT 9.225000  1.945000  9.555000 3.245000 ;
      RECT 9.295000  0.255000  9.485000 0.870000 ;
      RECT 9.655000  0.085000  9.985000 1.040000 ;
      RECT 9.725000  1.775000  9.985000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__a221oi_4
END LIBRARY
