* File: sky130_fd_sc_lp__a41o_2.pxi.spice
* Created: Wed Sep  2 09:29:01 2020
* 
x_PM_SKY130_FD_SC_LP__A41O_2%A_90_53# N_A_90_53#_M1002_s N_A_90_53#_M1003_d
+ N_A_90_53#_M1005_s N_A_90_53#_c_79_n N_A_90_53#_M1008_g N_A_90_53#_M1004_g
+ N_A_90_53#_c_81_n N_A_90_53#_M1011_g N_A_90_53#_M1013_g N_A_90_53#_c_82_n
+ N_A_90_53#_c_83_n N_A_90_53#_c_84_n N_A_90_53#_c_85_n N_A_90_53#_c_95_n
+ N_A_90_53#_c_96_n N_A_90_53#_c_97_n N_A_90_53#_c_86_n N_A_90_53#_c_87_n
+ N_A_90_53#_c_88_n N_A_90_53#_c_89_n N_A_90_53#_c_90_n
+ PM_SKY130_FD_SC_LP__A41O_2%A_90_53#
x_PM_SKY130_FD_SC_LP__A41O_2%B1 N_B1_M1002_g N_B1_M1005_g B1 N_B1_c_171_n
+ N_B1_c_172_n PM_SKY130_FD_SC_LP__A41O_2%B1
x_PM_SKY130_FD_SC_LP__A41O_2%A4 N_A4_M1001_g N_A4_M1006_g A4 N_A4_c_204_n
+ N_A4_c_205_n PM_SKY130_FD_SC_LP__A41O_2%A4
x_PM_SKY130_FD_SC_LP__A41O_2%A3 N_A3_M1007_g N_A3_M1012_g A3 N_A3_c_240_n
+ N_A3_c_241_n PM_SKY130_FD_SC_LP__A41O_2%A3
x_PM_SKY130_FD_SC_LP__A41O_2%A2 N_A2_M1009_g N_A2_M1000_g A2 A2 N_A2_c_277_n
+ PM_SKY130_FD_SC_LP__A41O_2%A2
x_PM_SKY130_FD_SC_LP__A41O_2%A1 N_A1_M1003_g N_A1_M1010_g A1 N_A1_c_312_n
+ N_A1_c_313_n PM_SKY130_FD_SC_LP__A41O_2%A1
x_PM_SKY130_FD_SC_LP__A41O_2%VPWR N_VPWR_M1004_d N_VPWR_M1013_d N_VPWR_M1001_d
+ N_VPWR_M1000_d N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n
+ N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n
+ VPWR N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_334_n N_VPWR_c_347_n
+ PM_SKY130_FD_SC_LP__A41O_2%VPWR
x_PM_SKY130_FD_SC_LP__A41O_2%X N_X_M1008_d N_X_M1004_s X X X X X X X
+ PM_SKY130_FD_SC_LP__A41O_2%X
x_PM_SKY130_FD_SC_LP__A41O_2%A_453_367# N_A_453_367#_M1005_d
+ N_A_453_367#_M1012_d N_A_453_367#_M1010_d N_A_453_367#_c_419_n
+ N_A_453_367#_c_442_n N_A_453_367#_c_421_n N_A_453_367#_c_427_n
+ N_A_453_367#_c_431_n N_A_453_367#_c_417_n N_A_453_367#_c_418_n
+ N_A_453_367#_c_428_n PM_SKY130_FD_SC_LP__A41O_2%A_453_367#
x_PM_SKY130_FD_SC_LP__A41O_2%VGND N_VGND_M1008_s N_VGND_M1011_s N_VGND_M1002_d
+ N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n
+ N_VGND_c_459_n VGND N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n
+ N_VGND_c_463_n PM_SKY130_FD_SC_LP__A41O_2%VGND
cc_1 VNB N_A_90_53#_c_79_n 0.0192049f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.345
cc_2 VNB N_A_90_53#_M1004_g 0.0127435f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_3 VNB N_A_90_53#_c_81_n 0.0389709f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.42
cc_4 VNB N_A_90_53#_c_82_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.42
cc_5 VNB N_A_90_53#_c_83_n 0.00744285f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.51
cc_6 VNB N_A_90_53#_c_84_n 0.0172692f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=0.42
cc_7 VNB N_A_90_53#_c_85_n 0.00623836f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=1.345
cc_8 VNB N_A_90_53#_c_86_n 0.0334151f $X=-0.19 $Y=-0.245 $X2=4.22 $Y2=1.08
cc_9 VNB N_A_90_53#_c_87_n 0.0288914f $X=-0.19 $Y=-0.245 $X2=4.385 $Y2=0.42
cc_10 VNB N_A_90_53#_c_88_n 0.00899941f $X=-0.19 $Y=-0.245 $X2=1.792 $Y2=1.08
cc_11 VNB N_A_90_53#_c_89_n 0.00553433f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=1.51
cc_12 VNB N_A_90_53#_c_90_n 0.0186192f $X=-0.19 $Y=-0.245 $X2=1.077 $Y2=1.345
cc_13 VNB N_B1_M1002_g 0.0300154f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.835
cc_14 VNB N_B1_c_171_n 0.0279984f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.815
cc_15 VNB N_B1_c_172_n 0.00328403f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.495
cc_16 VNB N_A4_M1006_g 0.0242456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A4_c_204_n 0.0262301f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.815
cc_18 VNB N_A4_c_205_n 0.00169879f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.495
cc_19 VNB N_A3_M1007_g 0.0242456f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.835
cc_20 VNB N_A3_c_240_n 0.0240969f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.815
cc_21 VNB N_A3_c_241_n 0.00357318f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.495
cc_22 VNB N_A2_M1009_g 0.0269114f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.835
cc_23 VNB A2 0.00462458f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.345
cc_24 VNB N_A2_c_277_n 0.0217423f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_25 VNB N_A1_M1003_g 0.0298742f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.835
cc_26 VNB N_A1_M1010_g 0.00138272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_c_312_n 0.0607015f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_28 VNB N_A1_c_313_n 0.0131744f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_29 VNB N_VPWR_c_334_n 0.203486f $X=-0.19 $Y=-0.245 $X2=1.077 $Y2=1.345
cc_30 VNB X 0.00717451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_454_n 0.0123082f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.345
cc_32 VNB N_VGND_c_455_n 0.0508265f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.815
cc_33 VNB N_VGND_c_456_n 0.0154949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_457_n 0.00599465f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.815
cc_35 VNB N_VGND_c_458_n 0.0250949f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.465
cc_36 VNB N_VGND_c_459_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.465
cc_37 VNB N_VGND_c_460_n 0.0164364f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.51
cc_38 VNB N_VGND_c_461_n 0.0681429f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=2.1
cc_39 VNB N_VGND_c_462_n 0.275768f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=2.91
cc_40 VNB N_VGND_c_463_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=4.385 $Y2=0.42
cc_41 VPB N_A_90_53#_M1004_g 0.0272005f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_42 VPB N_A_90_53#_c_81_n 0.00753942f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=1.42
cc_43 VPB N_A_90_53#_M1013_g 0.0226057f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_44 VPB N_A_90_53#_c_83_n 0.00691727f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=1.51
cc_45 VPB N_A_90_53#_c_95_n 0.00735195f $X=-0.19 $Y=1.655 $X2=1.75 $Y2=1.92
cc_46 VPB N_A_90_53#_c_96_n 0.00912238f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=2.1
cc_47 VPB N_A_90_53#_c_97_n 0.0157141f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=2.91
cc_48 VPB N_A_90_53#_c_89_n 0.00687345f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=1.51
cc_49 VPB N_B1_M1005_g 0.0226701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B1_c_171_n 0.0063819f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.815
cc_51 VPB N_B1_c_172_n 0.0047973f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.495
cc_52 VPB N_A4_M1001_g 0.0187338f $X=-0.19 $Y=1.655 $X2=1.85 $Y2=1.835
cc_53 VPB N_A4_c_204_n 0.0064469f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.815
cc_54 VPB N_A4_c_205_n 0.00257894f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.495
cc_55 VPB N_A3_M1012_g 0.0207713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A3_c_240_n 0.00624775f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.815
cc_57 VPB N_A3_c_241_n 0.00275689f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.495
cc_58 VPB N_A2_M1000_g 0.0203624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB A2 0.00499079f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.345
cc_60 VPB N_A2_c_277_n 0.00624794f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_61 VPB N_A1_M1010_g 0.0248773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A1_c_313_n 0.0121156f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_63 VPB N_VPWR_c_335_n 0.0122823f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.495
cc_64 VPB N_VPWR_c_336_n 0.0579608f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_65 VPB N_VPWR_c_337_n 0.022445f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=0.815
cc_66 VPB N_VPWR_c_338_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=1.505 $Y2=1.51
cc_67 VPB N_VPWR_c_339_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_340_n 0.0374261f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=0.42
cc_69 VPB N_VPWR_c_341_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_342_n 0.01926f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=1.345
cc_71 VPB N_VPWR_c_343_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.75 $Y2=1.675
cc_72 VPB N_VPWR_c_344_n 0.015372f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=2.91
cc_73 VPB N_VPWR_c_345_n 0.0203083f $X=-0.19 $Y=1.655 $X2=1.077 $Y2=1.42
cc_74 VPB N_VPWR_c_334_n 0.0731155f $X=-0.19 $Y=1.655 $X2=1.077 $Y2=1.345
cc_75 VPB N_VPWR_c_347_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB X 0.00456328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_453_367#_c_417_n 0.00785886f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=1.675
cc_78 VPB N_A_453_367#_c_418_n 0.0369431f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.465
cc_79 N_A_90_53#_c_85_n N_B1_M1002_g 0.00588467f $X=1.67 $Y=1.345 $X2=0 $Y2=0
cc_80 N_A_90_53#_c_86_n N_B1_M1002_g 0.0154097f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_81 N_A_90_53#_c_95_n N_B1_M1005_g 0.00512288f $X=1.75 $Y=1.92 $X2=0 $Y2=0
cc_82 N_A_90_53#_c_81_n N_B1_c_171_n 0.00355043f $X=0.88 $Y=1.42 $X2=0 $Y2=0
cc_83 N_A_90_53#_c_96_n N_B1_c_171_n 0.00286297f $X=1.945 $Y=2.1 $X2=0 $Y2=0
cc_84 N_A_90_53#_c_86_n N_B1_c_171_n 2.41424e-19 $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_85 N_A_90_53#_c_88_n N_B1_c_171_n 0.00370278f $X=1.792 $Y=1.08 $X2=0 $Y2=0
cc_86 N_A_90_53#_c_89_n N_B1_c_171_n 0.0042417f $X=1.67 $Y=1.51 $X2=0 $Y2=0
cc_87 N_A_90_53#_c_95_n N_B1_c_172_n 0.00586354f $X=1.75 $Y=1.92 $X2=0 $Y2=0
cc_88 N_A_90_53#_c_96_n N_B1_c_172_n 0.00510661f $X=1.945 $Y=2.1 $X2=0 $Y2=0
cc_89 N_A_90_53#_c_86_n N_B1_c_172_n 0.016021f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_90 N_A_90_53#_c_88_n N_B1_c_172_n 0.00609011f $X=1.792 $Y=1.08 $X2=0 $Y2=0
cc_91 N_A_90_53#_c_89_n N_B1_c_172_n 0.0276469f $X=1.67 $Y=1.51 $X2=0 $Y2=0
cc_92 N_A_90_53#_c_86_n N_A4_M1006_g 0.0151333f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_93 N_A_90_53#_c_86_n N_A4_c_204_n 0.00123623f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_94 N_A_90_53#_c_86_n N_A4_c_205_n 0.0235344f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_95 N_A_90_53#_c_86_n N_A3_M1007_g 0.0151473f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_96 N_A_90_53#_c_86_n N_A3_c_240_n 0.00249143f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_97 N_A_90_53#_c_86_n N_A3_c_241_n 0.0236976f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_98 N_A_90_53#_c_86_n N_A2_M1009_g 0.0161752f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_99 N_A_90_53#_c_87_n N_A2_M1009_g 0.00342706f $X=4.385 $Y=0.42 $X2=0 $Y2=0
cc_100 N_A_90_53#_c_86_n A2 0.0515643f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_101 N_A_90_53#_c_86_n N_A2_c_277_n 0.00443852f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_102 N_A_90_53#_c_86_n N_A1_M1003_g 0.0163323f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_103 N_A_90_53#_c_87_n N_A1_M1003_g 0.0175366f $X=4.385 $Y=0.42 $X2=0 $Y2=0
cc_104 N_A_90_53#_c_86_n N_A1_c_312_n 0.00970803f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_105 N_A_90_53#_c_86_n N_A1_c_313_n 0.0167876f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_106 N_A_90_53#_M1004_g N_VPWR_c_336_n 0.00757458f $X=0.525 $Y=2.465 $X2=0
+ $Y2=0
cc_107 N_A_90_53#_M1004_g N_VPWR_c_337_n 0.00112388f $X=0.525 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_90_53#_c_81_n N_VPWR_c_337_n 0.00553375f $X=0.88 $Y=1.42 $X2=0 $Y2=0
cc_109 N_A_90_53#_M1013_g N_VPWR_c_337_n 0.0222144f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_90_53#_c_83_n N_VPWR_c_337_n 0.0232149f $X=1.505 $Y=1.51 $X2=0 $Y2=0
cc_111 N_A_90_53#_c_95_n N_VPWR_c_337_n 0.00375739f $X=1.75 $Y=1.92 $X2=0 $Y2=0
cc_112 N_A_90_53#_c_96_n N_VPWR_c_337_n 0.00955412f $X=1.945 $Y=2.1 $X2=0 $Y2=0
cc_113 N_A_90_53#_c_97_n N_VPWR_c_337_n 0.0393049f $X=1.975 $Y=2.91 $X2=0 $Y2=0
cc_114 N_A_90_53#_c_97_n N_VPWR_c_340_n 0.0181659f $X=1.975 $Y=2.91 $X2=0 $Y2=0
cc_115 N_A_90_53#_M1004_g N_VPWR_c_344_n 0.00585385f $X=0.525 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_90_53#_M1013_g N_VPWR_c_344_n 0.00486043f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_90_53#_M1005_s N_VPWR_c_334_n 0.00336915f $X=1.85 $Y=1.835 $X2=0
+ $Y2=0
cc_118 N_A_90_53#_M1004_g N_VPWR_c_334_n 0.0116341f $X=0.525 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_A_90_53#_M1013_g N_VPWR_c_334_n 0.00835506f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_90_53#_c_97_n N_VPWR_c_334_n 0.0104192f $X=1.975 $Y=2.91 $X2=0 $Y2=0
cc_121 N_A_90_53#_c_79_n X 0.00340421f $X=0.525 $Y=1.345 $X2=0 $Y2=0
cc_122 N_A_90_53#_M1004_g X 0.00942991f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_90_53#_c_81_n X 0.0224696f $X=0.88 $Y=1.42 $X2=0 $Y2=0
cc_124 N_A_90_53#_c_83_n X 0.0240725f $X=1.505 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A_90_53#_c_85_n X 0.00430812f $X=1.67 $Y=1.345 $X2=0 $Y2=0
cc_126 N_A_90_53#_c_90_n X 0.00225116f $X=1.077 $Y=1.345 $X2=0 $Y2=0
cc_127 N_A_90_53#_c_86_n N_VGND_M1002_d 0.00308172f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_128 N_A_90_53#_c_79_n N_VGND_c_455_n 0.00725225f $X=0.525 $Y=1.345 $X2=0
+ $Y2=0
cc_129 N_A_90_53#_c_79_n N_VGND_c_456_n 5.15442e-19 $X=0.525 $Y=1.345 $X2=0
+ $Y2=0
cc_130 N_A_90_53#_c_81_n N_VGND_c_456_n 0.00553375f $X=0.88 $Y=1.42 $X2=0 $Y2=0
cc_131 N_A_90_53#_c_83_n N_VGND_c_456_n 0.0232149f $X=1.505 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A_90_53#_c_84_n N_VGND_c_456_n 0.0642696f $X=1.975 $Y=0.42 $X2=0 $Y2=0
cc_133 N_A_90_53#_c_85_n N_VGND_c_456_n 7.91056e-19 $X=1.67 $Y=1.345 $X2=0 $Y2=0
cc_134 N_A_90_53#_c_88_n N_VGND_c_456_n 0.0150383f $X=1.792 $Y=1.08 $X2=0 $Y2=0
cc_135 N_A_90_53#_c_90_n N_VGND_c_456_n 0.0169082f $X=1.077 $Y=1.345 $X2=0 $Y2=0
cc_136 N_A_90_53#_c_86_n N_VGND_c_457_n 0.022455f $X=4.22 $Y=1.08 $X2=0 $Y2=0
cc_137 N_A_90_53#_c_84_n N_VGND_c_458_n 0.0400304f $X=1.975 $Y=0.42 $X2=0 $Y2=0
cc_138 N_A_90_53#_c_79_n N_VGND_c_460_n 0.00559701f $X=0.525 $Y=1.345 $X2=0
+ $Y2=0
cc_139 N_A_90_53#_c_90_n N_VGND_c_460_n 0.00465077f $X=1.077 $Y=1.345 $X2=0
+ $Y2=0
cc_140 N_A_90_53#_c_87_n N_VGND_c_461_n 0.0210467f $X=4.385 $Y=0.42 $X2=0 $Y2=0
cc_141 N_A_90_53#_M1002_s N_VGND_c_462_n 0.00334057f $X=1.85 $Y=0.245 $X2=0
+ $Y2=0
cc_142 N_A_90_53#_M1003_d N_VGND_c_462_n 0.00212301f $X=4.245 $Y=0.245 $X2=0
+ $Y2=0
cc_143 N_A_90_53#_c_79_n N_VGND_c_462_n 0.00537853f $X=0.525 $Y=1.345 $X2=0
+ $Y2=0
cc_144 N_A_90_53#_c_84_n N_VGND_c_462_n 0.0222769f $X=1.975 $Y=0.42 $X2=0 $Y2=0
cc_145 N_A_90_53#_c_87_n N_VGND_c_462_n 0.0125689f $X=4.385 $Y=0.42 $X2=0 $Y2=0
cc_146 N_A_90_53#_c_90_n N_VGND_c_462_n 0.00451796f $X=1.077 $Y=1.345 $X2=0
+ $Y2=0
cc_147 N_A_90_53#_c_86_n A_561_49# 0.00366293f $X=4.22 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_90_53#_c_86_n A_633_49# 0.0106787f $X=4.22 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_90_53#_c_86_n A_741_49# 0.0106787f $X=4.22 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_150 N_B1_M1005_g N_A4_M1001_g 0.018713f $X=2.19 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B1_c_172_n N_A4_M1001_g 2.18895e-19 $X=2.1 $Y=1.51 $X2=0 $Y2=0
cc_152 N_B1_M1002_g N_A4_M1006_g 0.0181021f $X=2.19 $Y=0.665 $X2=0 $Y2=0
cc_153 N_B1_c_171_n N_A4_c_204_n 0.0206294f $X=2.1 $Y=1.51 $X2=0 $Y2=0
cc_154 N_B1_c_172_n N_A4_c_204_n 0.00184128f $X=2.1 $Y=1.51 $X2=0 $Y2=0
cc_155 N_B1_M1005_g N_A4_c_205_n 2.38927e-19 $X=2.19 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B1_c_171_n N_A4_c_205_n 3.80681e-19 $X=2.1 $Y=1.51 $X2=0 $Y2=0
cc_157 N_B1_c_172_n N_A4_c_205_n 0.0321181f $X=2.1 $Y=1.51 $X2=0 $Y2=0
cc_158 N_B1_M1005_g N_VPWR_c_338_n 0.00126699f $X=2.19 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B1_M1005_g N_VPWR_c_340_n 0.00585385f $X=2.19 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B1_M1005_g N_VPWR_c_334_n 0.0120903f $X=2.19 $Y=2.465 $X2=0 $Y2=0
cc_161 N_B1_M1002_g N_VGND_c_457_n 0.00312464f $X=2.19 $Y=0.665 $X2=0 $Y2=0
cc_162 N_B1_M1002_g N_VGND_c_458_n 0.00575161f $X=2.19 $Y=0.665 $X2=0 $Y2=0
cc_163 N_B1_M1002_g N_VGND_c_462_n 0.0121572f $X=2.19 $Y=0.665 $X2=0 $Y2=0
cc_164 N_A4_M1006_g N_A3_M1007_g 0.0497296f $X=2.73 $Y=0.665 $X2=0 $Y2=0
cc_165 N_A4_M1001_g N_A3_M1012_g 0.0320787f $X=2.62 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A4_c_205_n N_A3_M1012_g 2.46734e-19 $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A4_c_204_n N_A3_c_240_n 0.0497296f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_168 N_A4_c_205_n N_A3_c_240_n 3.80681e-19 $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A4_M1001_g N_A3_c_241_n 2.09427e-19 $X=2.62 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A4_c_204_n N_A3_c_241_n 0.00185954f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_171 N_A4_c_205_n N_A3_c_241_n 0.0323596f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A4_M1001_g N_VPWR_c_338_n 0.0139602f $X=2.62 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A4_M1001_g N_VPWR_c_340_n 0.00564095f $X=2.62 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A4_M1001_g N_VPWR_c_334_n 0.00950825f $X=2.62 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A4_c_204_n N_A_453_367#_c_419_n 2.02951e-19 $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A4_c_205_n N_A_453_367#_c_419_n 0.00244779f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A4_M1001_g N_A_453_367#_c_421_n 0.013307f $X=2.62 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A4_c_204_n N_A_453_367#_c_421_n 5.14933e-19 $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A4_c_205_n N_A_453_367#_c_421_n 0.0186539f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A4_M1006_g N_VGND_c_457_n 0.00312464f $X=2.73 $Y=0.665 $X2=0 $Y2=0
cc_181 N_A4_M1006_g N_VGND_c_461_n 0.00575161f $X=2.73 $Y=0.665 $X2=0 $Y2=0
cc_182 N_A4_M1006_g N_VGND_c_462_n 0.0107477f $X=2.73 $Y=0.665 $X2=0 $Y2=0
cc_183 N_A3_M1007_g N_A2_M1009_g 0.0443548f $X=3.09 $Y=0.665 $X2=0 $Y2=0
cc_184 N_A3_M1012_g N_A2_M1000_g 0.0278292f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A3_M1012_g A2 2.43457e-19 $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A3_c_240_n A2 0.00217937f $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_187 N_A3_c_241_n A2 0.0343715f $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A3_c_240_n N_A2_c_277_n 0.0205255f $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_189 N_A3_c_241_n N_A2_c_277_n 3.27415e-19 $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A3_M1012_g N_VPWR_c_338_n 0.0156124f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A3_M1012_g N_VPWR_c_339_n 9.95262e-19 $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A3_M1012_g N_VPWR_c_342_n 0.00564095f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A3_M1012_g N_VPWR_c_334_n 0.0100923f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A3_M1012_g N_A_453_367#_c_421_n 0.0165093f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A3_c_240_n N_A_453_367#_c_421_n 4.40054e-19 $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A3_c_241_n N_A_453_367#_c_421_n 0.0181364f $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A3_M1012_g N_A_453_367#_c_427_n 0.0131598f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A3_c_240_n N_A_453_367#_c_428_n 0.00196778f $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A3_c_241_n N_A_453_367#_c_428_n 0.00389035f $X=3.18 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A3_M1007_g N_VGND_c_461_n 0.00575161f $X=3.09 $Y=0.665 $X2=0 $Y2=0
cc_201 N_A3_M1007_g N_VGND_c_462_n 0.0109825f $X=3.09 $Y=0.665 $X2=0 $Y2=0
cc_202 N_A2_M1009_g N_A1_M1003_g 0.0407559f $X=3.63 $Y=0.665 $X2=0 $Y2=0
cc_203 N_A2_M1000_g N_A1_M1010_g 0.0376214f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_204 A2 N_A1_M1010_g 0.00421842f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_205 A2 N_A1_c_312_n 0.00987468f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_206 N_A2_c_277_n N_A1_c_312_n 0.0214326f $X=3.72 $Y=1.51 $X2=0 $Y2=0
cc_207 A2 N_A1_c_313_n 0.0329515f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_208 N_A2_M1000_g N_VPWR_c_338_n 9.8546e-19 $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A2_M1000_g N_VPWR_c_339_n 0.0165274f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A2_M1000_g N_VPWR_c_342_n 0.00486043f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A2_M1000_g N_VPWR_c_334_n 0.00885664f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A2_M1000_g N_A_453_367#_c_427_n 0.013109f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A2_M1000_g N_A_453_367#_c_431_n 0.0157149f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_214 A2 N_A_453_367#_c_431_n 0.0387169f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_215 N_A2_c_277_n N_A_453_367#_c_431_n 6.15792e-19 $X=3.72 $Y=1.51 $X2=0 $Y2=0
cc_216 A2 N_A_453_367#_c_428_n 0.0101206f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_217 N_A2_c_277_n N_A_453_367#_c_428_n 2.25908e-19 $X=3.72 $Y=1.51 $X2=0 $Y2=0
cc_218 N_A2_M1009_g N_VGND_c_461_n 0.00575161f $X=3.63 $Y=0.665 $X2=0 $Y2=0
cc_219 N_A2_M1009_g N_VGND_c_462_n 0.011406f $X=3.63 $Y=0.665 $X2=0 $Y2=0
cc_220 N_A1_M1010_g N_VPWR_c_339_n 0.0163574f $X=4.17 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A1_M1010_g N_VPWR_c_345_n 0.00486043f $X=4.17 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A1_M1010_g N_VPWR_c_334_n 0.00929712f $X=4.17 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A1_M1010_g N_A_453_367#_c_431_n 0.0146378f $X=4.17 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A1_c_312_n N_A_453_367#_c_417_n 0.00311076f $X=4.51 $Y=1.46 $X2=0 $Y2=0
cc_225 N_A1_c_313_n N_A_453_367#_c_417_n 0.0181076f $X=4.51 $Y=1.46 $X2=0 $Y2=0
cc_226 N_A1_M1003_g N_VGND_c_461_n 0.00539298f $X=4.17 $Y=0.665 $X2=0 $Y2=0
cc_227 N_A1_M1003_g N_VGND_c_462_n 0.0112898f $X=4.17 $Y=0.665 $X2=0 $Y2=0
cc_228 N_VPWR_c_334_n N_X_M1004_s 0.00392867f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_c_336_n X 0.0418332f $X=0.31 $Y=1.98 $X2=0 $Y2=0
cc_230 N_VPWR_c_344_n X 0.00857089f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_334_n X 0.00857956f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_232 N_VPWR_c_334_n N_A_453_367#_M1005_d 0.00432284f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_233 N_VPWR_c_334_n N_A_453_367#_M1012_d 0.0100514f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_334_n N_A_453_367#_M1010_d 0.00371702f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_340_n N_A_453_367#_c_442_n 0.0135169f $X=2.69 $Y=3.33 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_334_n N_A_453_367#_c_442_n 0.00847534f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_M1001_d N_A_453_367#_c_421_n 0.0085577f $X=2.695 $Y=1.835 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_338_n N_A_453_367#_c_421_n 0.0173521f $X=2.855 $Y=2.385 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_338_n N_A_453_367#_c_427_n 0.0479584f $X=2.855 $Y=2.385 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_339_n N_A_453_367#_c_427_n 0.0551387f $X=3.955 $Y=2.385 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_342_n N_A_453_367#_c_427_n 0.0230625f $X=3.79 $Y=3.33 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_334_n N_A_453_367#_c_427_n 0.0127519f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_VPWR_M1000_d N_A_453_367#_c_431_n 0.00351305f $X=3.815 $Y=1.835 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_339_n N_A_453_367#_c_431_n 0.0171443f $X=3.955 $Y=2.385 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_345_n N_A_453_367#_c_418_n 0.0178111f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_334_n N_A_453_367#_c_418_n 0.0100304f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_336_n N_VGND_c_455_n 0.011531f $X=0.31 $Y=1.98 $X2=0 $Y2=0
cc_248 N_VPWR_c_337_n N_VGND_c_456_n 5.07692e-19 $X=1.17 $Y=2.01 $X2=0 $Y2=0
cc_249 X N_VGND_c_455_n 0.0330999f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_250 X N_VGND_c_456_n 0.0319244f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_251 X N_VGND_c_460_n 0.00999534f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_252 X N_VGND_c_462_n 0.00855351f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_253 N_VGND_c_462_n A_561_49# 0.00899413f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
cc_254 N_VGND_c_462_n A_633_49# 0.0167034f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
cc_255 N_VGND_c_462_n A_741_49# 0.0167034f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
