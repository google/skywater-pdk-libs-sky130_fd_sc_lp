* File: sky130_fd_sc_lp__nor3_lp.pxi.spice
* Created: Fri Aug 28 10:55:51 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3_LP%C N_C_M1000_g N_C_c_52_n N_C_c_53_n N_C_M1002_g
+ N_C_c_58_n N_C_M1001_g N_C_c_55_n N_C_c_59_n C C N_C_c_57_n
+ PM_SKY130_FD_SC_LP__NOR3_LP%C
x_PM_SKY130_FD_SC_LP__NOR3_LP%B N_B_c_100_n N_B_M1006_g N_B_M1005_g N_B_c_101_n
+ N_B_M1003_g N_B_c_102_n N_B_c_103_n N_B_c_104_n N_B_c_109_n B B B B B
+ N_B_c_106_n PM_SKY130_FD_SC_LP__NOR3_LP%B
x_PM_SKY130_FD_SC_LP__NOR3_LP%A N_A_M1008_g N_A_c_162_n N_A_M1004_g N_A_M1007_g
+ N_A_c_163_n A A N_A_c_161_n PM_SKY130_FD_SC_LP__NOR3_LP%A
x_PM_SKY130_FD_SC_LP__NOR3_LP%Y N_Y_M1000_s N_Y_M1003_d N_Y_M1001_s N_Y_c_190_n
+ N_Y_c_191_n N_Y_c_192_n Y Y Y Y Y N_Y_c_194_n N_Y_c_196_n
+ PM_SKY130_FD_SC_LP__NOR3_LP%Y
x_PM_SKY130_FD_SC_LP__NOR3_LP%VPWR N_VPWR_M1004_d N_VPWR_c_244_n VPWR
+ N_VPWR_c_245_n N_VPWR_c_246_n N_VPWR_c_243_n N_VPWR_c_248_n
+ PM_SKY130_FD_SC_LP__NOR3_LP%VPWR
x_PM_SKY130_FD_SC_LP__NOR3_LP%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_c_264_n
+ N_VGND_c_265_n N_VGND_c_266_n VGND N_VGND_c_267_n N_VGND_c_268_n
+ N_VGND_c_269_n N_VGND_c_270_n PM_SKY130_FD_SC_LP__NOR3_LP%VGND
cc_1 VNB N_C_M1000_g 0.040069f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.495
cc_2 VNB N_C_c_52_n 0.0105634f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.25
cc_3 VNB N_C_c_53_n 0.0112215f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.25
cc_4 VNB N_C_M1002_g 0.0334464f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.495
cc_5 VNB N_C_c_55_n 0.0130831f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.25
cc_6 VNB C 0.00152213f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_7 VNB N_C_c_57_n 0.0267885f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.34
cc_8 VNB N_B_c_100_n 0.01389f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.175
cc_9 VNB N_B_c_101_n 0.0137713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_102_n 0.0214822f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.68
cc_11 VNB N_B_c_103_n 0.0156042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_104_n 0.0192294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB B 0.0118315f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.34
cc_14 VNB N_B_c_106_n 0.0130866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_M1008_g 0.0254837f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.495
cc_16 VNB N_A_M1007_g 0.0349485f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.545
cc_17 VNB A 0.0393902f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_18 VNB N_A_c_161_n 0.0731313f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.295
cc_19 VNB N_Y_c_190_n 0.0240181f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.545
cc_20 VNB N_Y_c_191_n 0.0214823f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.325
cc_21 VNB N_Y_c_192_n 0.0087472f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_22 VNB Y 0.0088017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_194_n 0.0489741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_243_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.34
cc_25 VNB N_VGND_c_264_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=0.495
cc_26 VNB N_VGND_c_265_n 0.015689f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.97
cc_27 VNB N_VGND_c_266_n 0.0253942f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.545
cc_28 VNB N_VGND_c_267_n 0.0365861f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_29 VNB N_VGND_c_268_n 0.0352342f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.34
cc_30 VNB N_VGND_c_269_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_270_n 0.224966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_C_c_58_n 0.0236431f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=1.97
cc_33 VPB N_C_c_59_n 0.0330459f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.68
cc_34 VPB C 0.00171029f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_35 VPB N_C_c_57_n 0.00195443f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.34
cc_36 VPB N_B_M1005_g 0.0262176f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=0.495
cc_37 VPB N_B_c_104_n 0.0018047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_B_c_109_n 0.0125316f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.34
cc_39 VPB B 0.00750996f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.34
cc_40 VPB N_A_c_162_n 0.031138f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.175
cc_41 VPB N_A_c_163_n 0.0166587f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.325
cc_42 VPB A 0.0258213f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_43 VPB N_A_c_161_n 0.0124588f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.295
cc_44 VPB Y 0.0285615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_Y_c_196_n 0.0837818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_244_n 0.0464658f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.25
cc_47 VPB N_VPWR_c_245_n 0.0686618f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.545
cc_48 VPB N_VPWR_c_246_n 0.0183725f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.34
cc_49 VPB N_VPWR_c_243_n 0.0798368f $X=-0.19 $Y=1.655 $X2=1.22 $Y2=1.34
cc_50 VPB N_VPWR_c_248_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 N_C_M1002_g N_B_c_100_n 0.0197172f $X=1.15 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_52 N_C_c_58_n N_B_M1005_g 0.0351035f $X=1.36 $Y=1.97 $X2=0 $Y2=0
cc_53 N_C_M1002_g N_B_c_103_n 0.00662647f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_54 N_C_c_55_n N_B_c_103_n 0.00745328f $X=1.22 $Y=1.25 $X2=0 $Y2=0
cc_55 N_C_c_59_n N_B_c_104_n 0.00745328f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_56 N_C_c_59_n N_B_c_109_n 0.0351035f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_57 N_C_c_55_n B 0.00529792f $X=1.22 $Y=1.25 $X2=0 $Y2=0
cc_58 N_C_c_59_n B 0.0141929f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_59 C B 0.0536046f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_60 C N_B_c_106_n 6.59086e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_61 N_C_c_57_n N_B_c_106_n 0.00745328f $X=1.22 $Y=1.34 $X2=0 $Y2=0
cc_62 N_C_M1000_g N_Y_c_190_n 0.01276f $X=0.79 $Y=0.495 $X2=0 $Y2=0
cc_63 N_C_M1002_g N_Y_c_190_n 0.00193397f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_64 N_C_M1000_g N_Y_c_191_n 0.00382866f $X=0.79 $Y=0.495 $X2=0 $Y2=0
cc_65 N_C_c_52_n N_Y_c_191_n 0.00101607f $X=1.055 $Y=1.25 $X2=0 $Y2=0
cc_66 N_C_M1002_g N_Y_c_191_n 0.011563f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_67 N_C_c_55_n N_Y_c_191_n 0.00109261f $X=1.22 $Y=1.25 $X2=0 $Y2=0
cc_68 C N_Y_c_191_n 0.0245017f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_69 N_C_c_59_n Y 0.00604189f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_70 C Y 0.021487f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_71 N_C_c_57_n Y 0.00700368f $X=1.22 $Y=1.34 $X2=0 $Y2=0
cc_72 N_C_M1000_g N_Y_c_194_n 0.0160312f $X=0.79 $Y=0.495 $X2=0 $Y2=0
cc_73 N_C_c_53_n N_Y_c_194_n 0.0106737f $X=0.865 $Y=1.25 $X2=0 $Y2=0
cc_74 N_C_M1002_g N_Y_c_194_n 0.00110545f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_75 C N_Y_c_194_n 0.0243784f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 N_C_c_57_n N_Y_c_194_n 0.00474375f $X=1.22 $Y=1.34 $X2=0 $Y2=0
cc_77 N_C_c_53_n N_Y_c_196_n 0.00602066f $X=0.865 $Y=1.25 $X2=0 $Y2=0
cc_78 N_C_c_58_n N_Y_c_196_n 0.01825f $X=1.36 $Y=1.97 $X2=0 $Y2=0
cc_79 N_C_c_59_n N_Y_c_196_n 0.00138993f $X=1.22 $Y=1.68 $X2=0 $Y2=0
cc_80 C N_Y_c_196_n 0.0172817f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_81 N_C_c_58_n N_VPWR_c_245_n 0.0085862f $X=1.36 $Y=1.97 $X2=0 $Y2=0
cc_82 N_C_c_58_n N_VPWR_c_243_n 0.0165862f $X=1.36 $Y=1.97 $X2=0 $Y2=0
cc_83 N_C_M1000_g N_VGND_c_264_n 0.00189426f $X=0.79 $Y=0.495 $X2=0 $Y2=0
cc_84 N_C_M1002_g N_VGND_c_264_n 0.0106455f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_85 N_C_M1000_g N_VGND_c_267_n 0.00502664f $X=0.79 $Y=0.495 $X2=0 $Y2=0
cc_86 N_C_M1002_g N_VGND_c_267_n 0.00445056f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_87 N_C_M1000_g N_VGND_c_270_n 0.00639688f $X=0.79 $Y=0.495 $X2=0 $Y2=0
cc_88 N_C_M1002_g N_VGND_c_270_n 0.0041956f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_89 N_B_c_101_n N_A_M1008_g 0.0169862f $X=1.94 $Y=0.78 $X2=0 $Y2=0
cc_90 N_B_c_103_n N_A_M1008_g 0.00785702f $X=1.89 $Y=1.18 $X2=0 $Y2=0
cc_91 N_B_M1005_g N_A_c_163_n 0.0483001f $X=1.85 $Y=2.545 $X2=0 $Y2=0
cc_92 N_B_c_104_n N_A_c_163_n 0.0175998f $X=1.89 $Y=1.685 $X2=0 $Y2=0
cc_93 N_B_c_103_n A 6.63751e-19 $X=1.89 $Y=1.18 $X2=0 $Y2=0
cc_94 B A 0.0405434f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B_c_106_n A 3.27326e-19 $X=1.89 $Y=1.345 $X2=0 $Y2=0
cc_96 B N_A_c_161_n 0.0198149f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B_c_106_n N_A_c_161_n 0.0175998f $X=1.89 $Y=1.345 $X2=0 $Y2=0
cc_98 N_B_c_102_n N_Y_c_191_n 0.0208196f $X=1.94 $Y=0.855 $X2=0 $Y2=0
cc_99 N_B_c_103_n N_Y_c_191_n 0.00495524f $X=1.89 $Y=1.18 $X2=0 $Y2=0
cc_100 B N_Y_c_191_n 0.0319023f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B_c_106_n N_Y_c_191_n 3.53153e-19 $X=1.89 $Y=1.345 $X2=0 $Y2=0
cc_102 N_B_c_100_n N_Y_c_192_n 0.00171214f $X=1.58 $Y=0.78 $X2=0 $Y2=0
cc_103 N_B_c_101_n N_Y_c_192_n 0.00975498f $X=1.94 $Y=0.78 $X2=0 $Y2=0
cc_104 N_B_c_102_n N_Y_c_192_n 0.00343296f $X=1.94 $Y=0.855 $X2=0 $Y2=0
cc_105 B N_Y_c_192_n 0.019925f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B_c_106_n N_Y_c_192_n 4.09568e-19 $X=1.89 $Y=1.345 $X2=0 $Y2=0
cc_107 N_B_M1005_g N_Y_c_196_n 0.00139793f $X=1.85 $Y=2.545 $X2=0 $Y2=0
cc_108 B N_Y_c_196_n 0.048165f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_109 B A_297_409# 0.0105574f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_110 B A_395_409# 0.00674313f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_111 N_B_M1005_g N_VPWR_c_244_n 0.00193455f $X=1.85 $Y=2.545 $X2=0 $Y2=0
cc_112 B N_VPWR_c_244_n 0.0248973f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B_M1005_g N_VPWR_c_245_n 0.00595064f $X=1.85 $Y=2.545 $X2=0 $Y2=0
cc_114 B N_VPWR_c_245_n 0.019793f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B_M1005_g N_VPWR_c_243_n 0.00772137f $X=1.85 $Y=2.545 $X2=0 $Y2=0
cc_116 B N_VPWR_c_243_n 0.0234398f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B_c_100_n N_VGND_c_264_n 0.0106389f $X=1.58 $Y=0.78 $X2=0 $Y2=0
cc_118 N_B_c_101_n N_VGND_c_264_n 0.00189367f $X=1.94 $Y=0.78 $X2=0 $Y2=0
cc_119 N_B_c_100_n N_VGND_c_268_n 0.00445056f $X=1.58 $Y=0.78 $X2=0 $Y2=0
cc_120 N_B_c_101_n N_VGND_c_268_n 0.00501274f $X=1.94 $Y=0.78 $X2=0 $Y2=0
cc_121 N_B_c_102_n N_VGND_c_268_n 5.84996e-19 $X=1.94 $Y=0.855 $X2=0 $Y2=0
cc_122 N_B_c_100_n N_VGND_c_270_n 0.0041956f $X=1.58 $Y=0.78 $X2=0 $Y2=0
cc_123 N_B_c_101_n N_VGND_c_270_n 0.00564643f $X=1.94 $Y=0.78 $X2=0 $Y2=0
cc_124 N_B_c_102_n N_VGND_c_270_n 7.94744e-19 $X=1.94 $Y=0.855 $X2=0 $Y2=0
cc_125 N_A_M1008_g N_Y_c_192_n 0.0167521f $X=2.37 $Y=0.495 $X2=0 $Y2=0
cc_126 N_A_M1007_g N_Y_c_192_n 0.00125398f $X=2.73 $Y=0.495 $X2=0 $Y2=0
cc_127 N_A_c_162_n N_VPWR_c_244_n 0.0220266f $X=2.42 $Y=2.04 $X2=0 $Y2=0
cc_128 A N_VPWR_c_244_n 0.0233028f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_129 N_A_c_161_n N_VPWR_c_244_n 0.00184748f $X=2.69 $Y=1.17 $X2=0 $Y2=0
cc_130 N_A_c_162_n N_VPWR_c_245_n 0.00802402f $X=2.42 $Y=2.04 $X2=0 $Y2=0
cc_131 N_A_c_162_n N_VPWR_c_243_n 0.0144019f $X=2.42 $Y=2.04 $X2=0 $Y2=0
cc_132 N_A_M1008_g N_VGND_c_266_n 0.00211129f $X=2.37 $Y=0.495 $X2=0 $Y2=0
cc_133 N_A_M1007_g N_VGND_c_266_n 0.0141573f $X=2.73 $Y=0.495 $X2=0 $Y2=0
cc_134 A N_VGND_c_266_n 0.0211412f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A_c_161_n N_VGND_c_266_n 0.00125242f $X=2.69 $Y=1.17 $X2=0 $Y2=0
cc_136 N_A_M1008_g N_VGND_c_268_n 0.00501274f $X=2.37 $Y=0.495 $X2=0 $Y2=0
cc_137 N_A_M1007_g N_VGND_c_268_n 0.00445056f $X=2.73 $Y=0.495 $X2=0 $Y2=0
cc_138 N_A_M1008_g N_VGND_c_270_n 0.00938368f $X=2.37 $Y=0.495 $X2=0 $Y2=0
cc_139 N_A_M1007_g N_VGND_c_270_n 0.00796275f $X=2.73 $Y=0.495 $X2=0 $Y2=0
cc_140 N_Y_c_196_n N_VPWR_c_245_n 0.0484708f $X=1.095 $Y=2.19 $X2=0 $Y2=0
cc_141 N_Y_c_196_n N_VPWR_c_243_n 0.0407141f $X=1.095 $Y=2.19 $X2=0 $Y2=0
cc_142 N_Y_c_190_n N_VGND_c_264_n 0.0127138f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_143 N_Y_c_191_n N_VGND_c_264_n 0.0200008f $X=1.99 $Y=0.91 $X2=0 $Y2=0
cc_144 N_Y_c_192_n N_VGND_c_264_n 0.0127434f $X=2.155 $Y=0.495 $X2=0 $Y2=0
cc_145 N_Y_c_192_n N_VGND_c_266_n 0.0154263f $X=2.155 $Y=0.495 $X2=0 $Y2=0
cc_146 N_Y_c_190_n N_VGND_c_267_n 0.0220321f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_147 N_Y_c_192_n N_VGND_c_268_n 0.0217716f $X=2.155 $Y=0.495 $X2=0 $Y2=0
cc_148 N_Y_c_190_n N_VGND_c_270_n 0.0125808f $X=0.575 $Y=0.495 $X2=0 $Y2=0
cc_149 N_Y_c_191_n N_VGND_c_270_n 0.0263778f $X=1.99 $Y=0.91 $X2=0 $Y2=0
cc_150 N_Y_c_192_n N_VGND_c_270_n 0.0124747f $X=2.155 $Y=0.495 $X2=0 $Y2=0
cc_151 N_Y_c_194_n N_VGND_c_270_n 0.00306138f $X=0.48 $Y=1.535 $X2=0 $Y2=0
