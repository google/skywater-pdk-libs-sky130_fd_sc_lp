* NGSPICE file created from sky130_fd_sc_lp__o21ba_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o21ba_0 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_499_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=3.78e+11p ps=3.48e+06u
M1001 VPWR a_80_225# X VPB phighvt w=640000u l=150000u
+  ad=6.581e+11p pd=6.12e+06u as=1.696e+11p ps=1.81e+06u
M1002 VGND a_80_225# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 a_557_487# A2 a_80_225# VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.792e+11p ps=1.84e+06u
M1004 a_499_47# a_258_397# a_80_225# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 a_80_225# a_258_397# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_258_397# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_258_397# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 VGND A2 a_499_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_557_487# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

