# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a2bb2oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.220000 1.405000 8.040000 1.755000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.210000 1.210000 8.965000 1.345000 ;
        RECT 8.210000 1.345000 9.560000 1.525000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.295000 1.350000 1.805000 1.555000 ;
        RECT 1.635000 1.555000 1.805000 1.665000 ;
        RECT 1.635000 1.665000 3.825000 1.835000 ;
        RECT 3.505000 1.200000 3.825000 1.665000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.315000 3.335000 1.485000 ;
        RECT 2.040000 1.200000 3.335000 1.315000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.050000 0.755000 4.545000 1.030000 ;
        RECT 3.995000 1.030000 4.165000 1.885000 ;
        RECT 3.995000 1.885000 4.770000 1.890000 ;
        RECT 3.995000 1.890000 5.545000 2.085000 ;
        RECT 4.310000 0.255000 4.545000 0.755000 ;
        RECT 4.345000 1.030000 4.545000 1.045000 ;
        RECT 4.345000 1.045000 5.700000 1.215000 ;
        RECT 4.355000 2.085000 4.685000 2.735000 ;
        RECT 5.215000 0.255000 5.405000 1.045000 ;
        RECT 5.215000 2.085000 5.545000 2.735000 ;
        RECT 5.355000 1.215000 5.700000 1.380000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.325000  1.725000  1.465000 1.895000 ;
      RECT 0.325000  1.895000  0.585000 3.075000 ;
      RECT 0.330000  0.085000  0.620000 1.095000 ;
      RECT 0.755000  2.065000  1.085000 3.245000 ;
      RECT 0.790000  0.255000  1.020000 1.010000 ;
      RECT 0.790000  1.010000  1.870000 1.180000 ;
      RECT 1.190000  0.085000  1.520000 0.840000 ;
      RECT 1.255000  1.895000  1.465000 2.015000 ;
      RECT 1.255000  2.015000  3.715000 2.185000 ;
      RECT 1.255000  2.185000  1.445000 3.075000 ;
      RECT 1.615000  2.355000  1.945000 3.245000 ;
      RECT 1.690000  0.255000  3.640000 0.585000 ;
      RECT 1.690000  0.585000  1.870000 1.010000 ;
      RECT 2.115000  2.185000  2.305000 3.075000 ;
      RECT 2.475000  2.355000  2.805000 3.245000 ;
      RECT 2.975000  2.185000  3.715000 2.245000 ;
      RECT 2.975000  2.245000  3.905000 2.255000 ;
      RECT 2.975000  2.255000  4.185000 2.415000 ;
      RECT 2.975000  2.415000  3.175000 3.075000 ;
      RECT 3.415000  2.585000  3.745000 3.245000 ;
      RECT 3.810000  0.085000  4.140000 0.585000 ;
      RECT 3.845000  2.415000  4.185000 2.425000 ;
      RECT 3.915000  2.425000  4.185000 2.905000 ;
      RECT 3.915000  2.905000  5.975000 3.075000 ;
      RECT 4.335000  1.385000  5.185000 1.550000 ;
      RECT 4.335000  1.550000  6.050000 1.715000 ;
      RECT 4.715000  0.085000  5.045000 0.865000 ;
      RECT 4.855000  2.255000  5.045000 2.905000 ;
      RECT 4.940000  1.715000  6.050000 1.720000 ;
      RECT 5.575000  0.085000  5.905000 0.875000 ;
      RECT 5.715000  1.890000  5.975000 2.905000 ;
      RECT 5.880000  1.065000  8.040000 1.235000 ;
      RECT 5.880000  1.235000  6.050000 1.550000 ;
      RECT 6.075000  0.255000  6.265000 1.065000 ;
      RECT 6.165000  1.930000  8.170000 2.100000 ;
      RECT 6.165000  2.100000  6.425000 3.075000 ;
      RECT 6.435000  0.085000  6.765000 0.895000 ;
      RECT 6.595000  2.270000  6.925000 3.245000 ;
      RECT 6.935000  0.255000  7.125000 1.040000 ;
      RECT 6.935000  1.040000  8.040000 1.065000 ;
      RECT 7.095000  2.100000  7.285000 3.075000 ;
      RECT 7.295000  0.085000  8.135000 0.700000 ;
      RECT 7.295000  0.700000  7.625000 0.870000 ;
      RECT 7.455000  2.270000  7.785000 3.245000 ;
      RECT 7.870000  0.870000  9.365000 1.005000 ;
      RECT 7.870000  1.005000  9.935000 1.040000 ;
      RECT 7.955000  2.100000  8.170000 2.905000 ;
      RECT 7.955000  2.905000  9.935000 3.075000 ;
      RECT 8.305000  0.255000  8.505000 0.870000 ;
      RECT 8.340000  1.695000  9.935000 1.875000 ;
      RECT 8.340000  1.875000  8.615000 2.735000 ;
      RECT 8.675000  0.085000  9.005000 0.700000 ;
      RECT 8.785000  2.045000  9.045000 2.905000 ;
      RECT 9.165000  1.040000  9.935000 1.175000 ;
      RECT 9.175000  0.255000  9.365000 0.870000 ;
      RECT 9.215000  1.875000  9.475000 2.735000 ;
      RECT 9.535000  0.085000  9.865000 0.835000 ;
      RECT 9.645000  2.045000  9.935000 2.905000 ;
      RECT 9.730000  1.175000  9.935000 1.695000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__a2bb2oi_4
END LIBRARY
