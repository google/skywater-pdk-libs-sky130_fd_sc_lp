* NGSPICE file created from sky130_fd_sc_lp__ebufn_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__ebufn_4 A TE_B VGND VNB VPB VPWR Z
M1000 Z a_84_21# a_27_47# VNB nshort w=840000u l=150000u
+  ad=5.292e+11p pd=4.62e+06u as=1.2432e+12p ps=1.136e+07u
M1001 Z a_84_21# a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.938e+11p pd=6.3e+06u as=1.953e+12p ps=1.57e+07u
M1002 VPWR TE_B a_456_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.5498e+12p pd=1.002e+07u as=5.185e+11p ps=3.42e+06u
M1003 a_27_47# a_84_21# Z VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Z a_84_21# a_27_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_84_21# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1006 a_27_367# a_84_21# Z VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_367# TE_B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_456_21# a_27_47# VNB nshort w=840000u l=150000u
+  ad=8.232e+11p pd=7e+06u as=0p ps=0u
M1009 VPWR TE_B a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_456_21# a_27_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Z a_84_21# a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND TE_B a_456_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1013 a_27_47# a_456_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_47# a_456_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_367# a_84_21# Z VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR TE_B a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_367# TE_B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_47# a_84_21# Z VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_84_21# A VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
.ends

