* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4bb_m A_N B_N C D VGND VNB VPB VPWR Y
X0 VPWR a_27_151# Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_427_151# a_469_125# Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_151# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_319_151# a_27_151# a_427_151# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_151# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 Y a_469_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND A_N a_469_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR A_N a_469_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND D a_247_151# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_247_151# C a_319_151# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
