* File: sky130_fd_sc_lp__mux2_1.spice
* Created: Wed Sep  2 10:00:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2_1.pex.spice"
.subckt sky130_fd_sc_lp__mux2_1  VNB VPB S A1 A0 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_105_22#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2156 AS=0.2226 PD=1.79333 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1007 A_266_132# N_S_M1007_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0672
+ AS=0.1078 PD=0.74 PS=0.896667 NRD=30 NRS=65.712 M=1 R=2.8 SA=75000.8
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_105_22#_M1001_d N_A1_M1001_g A_266_132# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75001.3
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1010 A_446_132# N_A0_M1010_g N_A_105_22#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_488_106#_M1008_g A_446_132# VNB NSHORT L=0.15 W=0.42
+ AD=0.1953 AS=0.0441 PD=1.35 PS=0.63 NRD=74.28 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_488_106#_M1003_d N_S_M1003_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1953 PD=1.41 PS=1.35 NRD=5.712 NRS=0 M=1 R=2.8 SA=75003.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_105_22#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.360675 AS=0.3339 PD=2.8125 PS=3.05 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1004 A_288_434# N_S_M1004_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.120225 PD=0.63 PS=0.9375 NRD=23.443 NRS=100.844 M=1 R=2.8 SA=75001
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1005 N_A_105_22#_M1005_d N_A0_M1005_g A_288_434# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1344 AS=0.0441 PD=1.06 PS=0.63 NRD=114.91 NRS=23.443 M=1 R=2.8 SA=75001.3
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1009 A_518_434# N_A1_M1009_g N_A_105_22#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1344 PD=0.81 PS=1.06 NRD=65.6601 NRS=53.9386 M=1 R=2.8
+ SA=75002.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_488_106#_M1000_g A_518_434# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=37.5088 NRS=65.6601 M=1 R=2.8
+ SA=75002.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_A_488_106#_M1011_d N_S_M1011_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=14.0658 M=1 R=2.8 SA=75003.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__mux2_1.pxi.spice"
*
.ends
*
*
