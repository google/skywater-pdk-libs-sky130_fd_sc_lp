* File: sky130_fd_sc_lp__a221oi_4.pex.spice
* Created: Wed Sep  2 09:22:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221OI_4%C1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 33 39 54
c88 24 0 2.45799e-20 $X=2.055 $Y=2.465
r89 52 54 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.09 $Y=1.35
+ $X2=2.225 $Y2=1.35
r90 50 52 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.055 $Y=1.35
+ $X2=2.09 $Y2=1.35
r91 49 50 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.795 $Y=1.35
+ $X2=2.055 $Y2=1.35
r92 48 49 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.625 $Y=1.35
+ $X2=1.795 $Y2=1.35
r93 47 48 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.365 $Y=1.35
+ $X2=1.625 $Y2=1.35
r94 46 47 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.195 $Y=1.35
+ $X2=1.365 $Y2=1.35
r95 45 46 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=0.935 $Y=1.35
+ $X2=1.195 $Y2=1.35
r96 44 45 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.765 $Y=1.35
+ $X2=0.935 $Y2=1.35
r97 41 42 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.39
+ $Y=1.35 $X2=0.39 $Y2=1.35
r98 39 44 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.69 $Y=1.35
+ $X2=0.765 $Y2=1.35
r99 39 41 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=0.69 $Y=1.35 $X2=0.39
+ $Y2=1.35
r100 33 52 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.09
+ $Y=1.35 $X2=2.09 $Y2=1.35
r101 32 33 21.0001 $w=2.23e-07 $l=4.1e-07 $layer=LI1_cond $X=1.68 $Y=1.322
+ $X2=2.09 $Y2=1.322
r102 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.322
+ $X2=1.68 $Y2=1.322
r103 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.322
+ $X2=1.2 $Y2=1.322
r104 30 42 16.9025 $w=2.23e-07 $l=3.3e-07 $layer=LI1_cond $X=0.72 $Y=1.322
+ $X2=0.39 $Y2=1.322
r105 29 42 7.68295 $w=2.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=1.322
+ $X2=0.39 $Y2=1.322
r106 26 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.185
+ $X2=2.225 $Y2=1.35
r107 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.225 $Y=1.185
+ $X2=2.225 $Y2=0.655
r108 22 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.055 $Y=1.515
+ $X2=2.055 $Y2=1.35
r109 22 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.055 $Y=1.515
+ $X2=2.055 $Y2=2.465
r110 19 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.185
+ $X2=1.795 $Y2=1.35
r111 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.795 $Y=1.185
+ $X2=1.795 $Y2=0.655
r112 15 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.515
+ $X2=1.625 $Y2=1.35
r113 15 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.625 $Y=1.515
+ $X2=1.625 $Y2=2.465
r114 12 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.185
+ $X2=1.365 $Y2=1.35
r115 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.365 $Y=1.185
+ $X2=1.365 $Y2=0.655
r116 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.515
+ $X2=1.195 $Y2=1.35
r117 8 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.195 $Y=1.515
+ $X2=1.195 $Y2=2.465
r118 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.185
+ $X2=0.935 $Y2=1.35
r119 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=1.185
+ $X2=0.935 $Y2=0.655
r120 1 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.765 $Y=1.515
+ $X2=0.765 $Y2=1.35
r121 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.765 $Y=1.515
+ $X2=0.765 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%B2 3 7 11 15 19 23 27 31 33 38 39 40 41 46
+ 57 60 61 70
c135 60 0 1.5135e-19 $X=6.035 $Y=1.51
c136 40 0 1.38485e-19 $X=5.85 $Y=2.015
c137 39 0 3.74771e-20 $X=3.73 $Y=1.93
c138 38 0 1.48878e-19 $X=3.73 $Y=1.625
c139 33 0 2.45799e-20 $X=3.645 $Y=1.525
c140 31 0 1.1786e-19 $X=6.085 $Y=0.655
r141 70 71 1.57788 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=6.025 $Y=1.665
+ $X2=6.025 $Y2=1.675
r142 60 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.035 $Y=1.51
+ $X2=6.035 $Y2=1.675
r143 60 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.035 $Y=1.51
+ $X2=6.035 $Y2=1.345
r144 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.035
+ $Y=1.51 $X2=6.035 $Y2=1.51
r145 54 55 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.435 $Y=1.51
+ $X2=3.515 $Y2=1.51
r146 53 54 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.085 $Y=1.51
+ $X2=3.435 $Y2=1.51
r147 52 53 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.005 $Y=1.51
+ $X2=3.085 $Y2=1.51
r148 46 70 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=6.025 $Y=1.627
+ $X2=6.025 $Y2=1.665
r149 46 61 3.85245 $w=3.48e-07 $l=1.17e-07 $layer=LI1_cond $X=6.025 $Y=1.627
+ $X2=6.025 $Y2=1.51
r150 46 71 1.81448 $w=2.33e-07 $l=3.7e-08 $layer=LI1_cond $X=5.967 $Y=1.712
+ $X2=5.967 $Y2=1.675
r151 45 46 10.6907 $w=2.33e-07 $l=2.18e-07 $layer=LI1_cond $X=5.967 $Y=1.93
+ $X2=5.967 $Y2=1.712
r152 44 57 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.65 $Y=1.51
+ $X2=3.865 $Y2=1.51
r153 44 55 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.65 $Y=1.51
+ $X2=3.515 $Y2=1.51
r154 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.65
+ $Y=1.51 $X2=3.65 $Y2=1.51
r155 40 45 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=5.85 $Y=2.015
+ $X2=5.967 $Y2=1.93
r156 40 41 132.765 $w=1.68e-07 $l=2.035e-06 $layer=LI1_cond $X=5.85 $Y=2.015
+ $X2=3.815 $Y2=2.015
r157 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.73 $Y=1.93
+ $X2=3.815 $Y2=2.015
r158 38 43 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.73 $Y=1.625 $X2=3.73
+ $Y2=1.525
r159 38 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.73 $Y=1.625
+ $X2=3.73 $Y2=1.93
r160 36 52 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.97 $Y=1.51
+ $X2=3.005 $Y2=1.51
r161 36 49 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.97 $Y=1.51
+ $X2=2.655 $Y2=1.51
r162 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.97
+ $Y=1.51 $X2=2.97 $Y2=1.51
r163 33 43 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=1.525
+ $X2=3.73 $Y2=1.525
r164 33 35 37.4318 $w=1.98e-07 $l=6.75e-07 $layer=LI1_cond $X=3.645 $Y=1.525
+ $X2=2.97 $Y2=1.525
r165 31 62 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.085 $Y=0.655
+ $X2=6.085 $Y2=1.345
r166 27 63 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.015 $Y=2.465
+ $X2=6.015 $Y2=1.675
r167 21 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.865 $Y=1.675
+ $X2=3.865 $Y2=1.51
r168 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.865 $Y=1.675
+ $X2=3.865 $Y2=2.465
r169 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.345
+ $X2=3.515 $Y2=1.51
r170 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.515 $Y=1.345
+ $X2=3.515 $Y2=0.655
r171 13 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.435 $Y=1.675
+ $X2=3.435 $Y2=1.51
r172 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.435 $Y=1.675
+ $X2=3.435 $Y2=2.465
r173 9 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.345
+ $X2=3.085 $Y2=1.51
r174 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.085 $Y=1.345
+ $X2=3.085 $Y2=0.655
r175 5 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.005 $Y=1.675
+ $X2=3.005 $Y2=1.51
r176 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.005 $Y=1.675
+ $X2=3.005 $Y2=2.465
r177 1 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.345
+ $X2=2.655 $Y2=1.51
r178 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.655 $Y=1.345
+ $X2=2.655 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 53
c74 53 0 1.86355e-19 $X=5.515 $Y=1.51
r75 53 54 10.5109 $w=3.21e-07 $l=7e-08 $layer=POLY_cond $X=5.515 $Y=1.51
+ $X2=5.585 $Y2=1.51
r76 51 53 27.028 $w=3.21e-07 $l=1.8e-07 $layer=POLY_cond $X=5.335 $Y=1.51
+ $X2=5.515 $Y2=1.51
r77 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.335
+ $Y=1.51 $X2=5.335 $Y2=1.51
r78 49 51 27.028 $w=3.21e-07 $l=1.8e-07 $layer=POLY_cond $X=5.155 $Y=1.51
+ $X2=5.335 $Y2=1.51
r79 48 49 10.5109 $w=3.21e-07 $l=7e-08 $layer=POLY_cond $X=5.085 $Y=1.51
+ $X2=5.155 $Y2=1.51
r80 47 48 54.0561 $w=3.21e-07 $l=3.6e-07 $layer=POLY_cond $X=4.725 $Y=1.51
+ $X2=5.085 $Y2=1.51
r81 46 47 10.5109 $w=3.21e-07 $l=7e-08 $layer=POLY_cond $X=4.655 $Y=1.51
+ $X2=4.725 $Y2=1.51
r82 44 46 51.053 $w=3.21e-07 $l=3.4e-07 $layer=POLY_cond $X=4.315 $Y=1.51
+ $X2=4.655 $Y2=1.51
r83 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.315
+ $Y=1.51 $X2=4.315 $Y2=1.51
r84 42 44 3.00312 $w=3.21e-07 $l=2e-08 $layer=POLY_cond $X=4.295 $Y=1.51
+ $X2=4.315 $Y2=1.51
r85 41 42 10.5109 $w=3.21e-07 $l=7e-08 $layer=POLY_cond $X=4.225 $Y=1.51
+ $X2=4.295 $Y2=1.51
r86 36 52 5.26425 $w=4.03e-07 $l=1.85e-07 $layer=LI1_cond $X=5.52 $Y=1.557
+ $X2=5.335 $Y2=1.557
r87 35 52 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=5.04 $Y=1.557
+ $X2=5.335 $Y2=1.557
r88 34 35 13.6586 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.557
+ $X2=5.04 $Y2=1.557
r89 34 45 6.97157 $w=4.03e-07 $l=2.45e-07 $layer=LI1_cond $X=4.56 $Y=1.557
+ $X2=4.315 $Y2=1.557
r90 33 45 6.68702 $w=4.03e-07 $l=2.35e-07 $layer=LI1_cond $X=4.08 $Y=1.557
+ $X2=4.315 $Y2=1.557
r91 29 54 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=1.675
+ $X2=5.585 $Y2=1.51
r92 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.585 $Y=1.675
+ $X2=5.585 $Y2=2.465
r93 25 53 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.515 $Y=1.345
+ $X2=5.515 $Y2=1.51
r94 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.515 $Y=1.345
+ $X2=5.515 $Y2=0.655
r95 21 49 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.675
+ $X2=5.155 $Y2=1.51
r96 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.155 $Y=1.675
+ $X2=5.155 $Y2=2.465
r97 17 48 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.085 $Y=1.345
+ $X2=5.085 $Y2=1.51
r98 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.085 $Y=1.345
+ $X2=5.085 $Y2=0.655
r99 13 47 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.725 $Y=1.675
+ $X2=4.725 $Y2=1.51
r100 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.725 $Y=1.675
+ $X2=4.725 $Y2=2.465
r101 9 46 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=1.345
+ $X2=4.655 $Y2=1.51
r102 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.655 $Y=1.345
+ $X2=4.655 $Y2=0.655
r103 5 42 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.675
+ $X2=4.295 $Y2=1.51
r104 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.295 $Y=1.675
+ $X2=4.295 $Y2=2.465
r105 1 41 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.225 $Y=1.345
+ $X2=4.225 $Y2=1.51
r106 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.225 $Y=1.345
+ $X2=4.225 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%A2 3 7 9 11 14 16 18 21 23 25 28 30 32 33
+ 35 36 40 41 42 43 60
c125 35 0 1.0586e-19 $X=6.575 $Y=1.51
c126 32 0 3.31495e-20 $X=8.365 $Y=1.435
c127 3 0 1.38485e-19 $X=6.565 $Y=2.465
r128 58 60 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=9.605 $Y=1.35
+ $X2=9.785 $Y2=1.35
r129 57 58 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=9.175 $Y=1.35
+ $X2=9.605 $Y2=1.35
r130 55 57 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=8.765 $Y=1.35
+ $X2=9.175 $Y2=1.35
r131 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.765
+ $Y=1.35 $X2=8.765 $Y2=1.35
r132 52 55 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.745 $Y=1.35
+ $X2=8.765 $Y2=1.35
r133 43 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.785
+ $Y=1.35 $X2=9.785 $Y2=1.35
r134 42 43 21.7684 $w=2.23e-07 $l=4.25e-07 $layer=LI1_cond $X=9.36 $Y=1.322
+ $X2=9.785 $Y2=1.322
r135 41 42 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.322
+ $X2=9.36 $Y2=1.322
r136 41 56 5.89026 $w=2.23e-07 $l=1.15e-07 $layer=LI1_cond $X=8.88 $Y=1.322
+ $X2=8.765 $Y2=1.322
r137 40 56 10.2861 $w=3.93e-07 $l=2.8e-07 $layer=LI1_cond $X=8.485 $Y=1.322
+ $X2=8.765 $Y2=1.322
r138 36 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.575 $Y=1.51
+ $X2=6.575 $Y2=1.675
r139 36 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.575 $Y=1.51
+ $X2=6.575 $Y2=1.345
r140 35 38 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=6.535 $Y=1.51
+ $X2=6.535 $Y2=1.7
r141 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.575
+ $Y=1.51 $X2=6.575 $Y2=1.51
r142 32 40 3.31033 $w=2.4e-07 $l=1.13e-07 $layer=LI1_cond $X=8.365 $Y=1.435
+ $X2=8.365 $Y2=1.322
r143 32 33 8.64332 $w=2.38e-07 $l=1.8e-07 $layer=LI1_cond $X=8.365 $Y=1.435
+ $X2=8.365 $Y2=1.615
r144 31 38 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=1.7
+ $X2=6.535 $Y2=1.7
r145 30 33 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=8.245 $Y=1.7
+ $X2=8.365 $Y2=1.615
r146 30 31 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=8.245 $Y=1.7
+ $X2=6.66 $Y2=1.7
r147 26 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.515
+ $X2=9.605 $Y2=1.35
r148 26 28 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.605 $Y=1.515
+ $X2=9.605 $Y2=2.465
r149 23 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.185
+ $X2=9.605 $Y2=1.35
r150 23 25 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.605 $Y=1.185
+ $X2=9.605 $Y2=0.655
r151 19 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.175 $Y=1.515
+ $X2=9.175 $Y2=1.35
r152 19 21 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.175 $Y=1.515
+ $X2=9.175 $Y2=2.465
r153 16 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.175 $Y=1.185
+ $X2=9.175 $Y2=1.35
r154 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.175 $Y=1.185
+ $X2=9.175 $Y2=0.655
r155 12 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.745 $Y=1.515
+ $X2=8.745 $Y2=1.35
r156 12 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.745 $Y=1.515
+ $X2=8.745 $Y2=2.465
r157 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.745 $Y=1.185
+ $X2=8.745 $Y2=1.35
r158 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.745 $Y=1.185
+ $X2=8.745 $Y2=0.655
r159 7 50 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.595 $Y=0.655
+ $X2=6.595 $Y2=1.345
r160 3 51 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.565 $Y=2.465
+ $X2=6.565 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%A1 1 3 6 8 10 13 15 17 18 20 21 23 25 27 28
+ 30 31 32 33 45
c85 45 0 3.31495e-20 $X=7.885 $Y=1.455
c86 23 0 1.59281e-19 $X=8.24 $Y=1.65
c87 21 0 5.71875e-20 $X=8.24 $Y=1.26
c88 6 0 1.0586e-19 $X=7.025 $Y=2.465
r89 43 45 12.0166 $w=3.61e-07 $l=9e-08 $layer=POLY_cond $X=7.795 $Y=1.455
+ $X2=7.885 $Y2=1.455
r90 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.795
+ $Y=1.35 $X2=7.795 $Y2=1.35
r91 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.115
+ $Y=1.35 $X2=7.115 $Y2=1.35
r92 33 44 6.13002 $w=2.33e-07 $l=1.25e-07 $layer=LI1_cond $X=7.92 $Y=1.317
+ $X2=7.795 $Y2=1.317
r93 32 44 17.4092 $w=2.33e-07 $l=3.55e-07 $layer=LI1_cond $X=7.44 $Y=1.317
+ $X2=7.795 $Y2=1.317
r94 32 40 15.938 $w=2.33e-07 $l=3.25e-07 $layer=LI1_cond $X=7.44 $Y=1.317
+ $X2=7.115 $Y2=1.317
r95 31 40 7.60122 $w=2.33e-07 $l=1.55e-07 $layer=LI1_cond $X=6.96 $Y=1.317
+ $X2=7.115 $Y2=1.317
r96 28 30 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.315 $Y=1.725
+ $X2=8.315 $Y2=2.465
r97 25 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.315 $Y=1.185
+ $X2=8.315 $Y2=0.655
r98 24 45 20.3347 $w=1.8e-07 $l=2.29456e-07 $layer=POLY_cond $X=7.96 $Y=1.65
+ $X2=7.885 $Y2=1.455
r99 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.24 $Y=1.65
+ $X2=8.315 $Y2=1.725
r100 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.24 $Y=1.65
+ $X2=7.96 $Y2=1.65
r101 22 45 20.3347 $w=1.8e-07 $l=2.29456e-07 $layer=POLY_cond $X=7.96 $Y=1.26
+ $X2=7.885 $Y2=1.455
r102 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.24 $Y=1.26
+ $X2=8.315 $Y2=1.185
r103 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.24 $Y=1.26
+ $X2=7.96 $Y2=1.26
r104 18 45 23.3725 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.885 $Y=1.725
+ $X2=7.885 $Y2=1.455
r105 18 20 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.885 $Y=1.725
+ $X2=7.885 $Y2=2.465
r106 15 45 23.3725 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.885 $Y=1.185
+ $X2=7.885 $Y2=1.455
r107 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.885 $Y=1.185
+ $X2=7.885 $Y2=0.655
r108 11 43 45.3961 $w=3.61e-07 $l=3.4e-07 $layer=POLY_cond $X=7.455 $Y=1.455
+ $X2=7.795 $Y2=1.455
r109 11 39 45.3961 $w=3.61e-07 $l=3.4e-07 $layer=POLY_cond $X=7.455 $Y=1.455
+ $X2=7.115 $Y2=1.455
r110 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.455 $Y=1.515
+ $X2=7.455 $Y2=2.465
r111 8 11 23.3725 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.455 $Y=1.185
+ $X2=7.455 $Y2=1.455
r112 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.455 $Y=1.185
+ $X2=7.455 $Y2=0.655
r113 4 39 12.0166 $w=3.61e-07 $l=9e-08 $layer=POLY_cond $X=7.025 $Y=1.455
+ $X2=7.115 $Y2=1.455
r114 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.025 $Y=1.515
+ $X2=7.025 $Y2=2.465
r115 1 4 23.3725 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=1.455
r116 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%A_85_367# 1 2 3 4 5 6 7 22 24 26 30 34 36
+ 37 38 41 48 52 58
c77 48 0 1.5135e-19 $X=5.8 $Y=2.435
r78 60 61 4.4265 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=2.03 $X2=3.19
+ $Y2=2.115
r79 58 60 2.98782 $w=2.68e-07 $l=7e-08 $layer=LI1_cond $X=3.19 $Y=1.96 $X2=3.19
+ $Y2=2.03
r80 46 48 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.94 $Y=2.435
+ $X2=5.8 $Y2=2.435
r81 44 46 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.08 $Y=2.435
+ $X2=4.94 $Y2=2.435
r82 42 63 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=3.325 $Y=2.435
+ $X2=3.225 $Y2=2.435
r83 42 44 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=3.325 $Y=2.435
+ $X2=4.08 $Y2=2.435
r84 41 63 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=2.27
+ $X2=3.225 $Y2=2.435
r85 41 61 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=3.225 $Y=2.27
+ $X2=3.225 $Y2=2.115
r86 39 54 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.435 $Y=2.03
+ $X2=2.305 $Y2=2.03
r87 38 60 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.055 $Y=2.03
+ $X2=3.19 $Y2=2.03
r88 38 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.055 $Y=2.03
+ $X2=2.435 $Y2=2.03
r89 37 56 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=2.905
+ $X2=2.305 $Y2=2.99
r90 36 54 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=2.115
+ $X2=2.305 $Y2=2.03
r91 36 37 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=2.305 $Y=2.115
+ $X2=2.305 $Y2=2.905
r92 35 52 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.505 $Y=2.99
+ $X2=1.41 $Y2=2.99
r93 34 56 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.175 $Y=2.99
+ $X2=2.305 $Y2=2.99
r94 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.175 $Y=2.99
+ $X2=1.505 $Y2=2.99
r95 30 33 45.5311 $w=1.88e-07 $l=7.8e-07 $layer=LI1_cond $X=1.41 $Y=2.11
+ $X2=1.41 $Y2=2.89
r96 28 52 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=2.905
+ $X2=1.41 $Y2=2.99
r97 28 33 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=1.41 $Y=2.905
+ $X2=1.41 $Y2=2.89
r98 27 51 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.645 $Y=2.99
+ $X2=0.515 $Y2=2.99
r99 26 52 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.315 $Y=2.99
+ $X2=1.41 $Y2=2.99
r100 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.315 $Y=2.99
+ $X2=0.645 $Y2=2.99
r101 22 51 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.515 $Y=2.905
+ $X2=0.515 $Y2=2.99
r102 22 24 41.0004 $w=2.58e-07 $l=9.25e-07 $layer=LI1_cond $X=0.515 $Y=2.905
+ $X2=0.515 $Y2=1.98
r103 7 48 600 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=1 $X=5.66
+ $Y=1.835 $X2=5.8 $Y2=2.435
r104 6 46 600 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=1.835 $X2=4.94 $Y2=2.435
r105 5 44 600 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=1.835 $X2=4.08 $Y2=2.435
r106 4 63 600 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.835 $X2=3.22 $Y2=2.435
r107 4 58 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.835 $X2=3.22 $Y2=1.96
r108 3 56 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.835 $X2=2.27 $Y2=2.91
r109 3 54 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.13
+ $Y=1.835 $X2=2.27 $Y2=2.11
r110 2 33 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=1.27
+ $Y=1.835 $X2=1.41 $Y2=2.89
r111 2 30 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.27
+ $Y=1.835 $X2=1.41 $Y2=2.11
r112 1 51 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.425
+ $Y=1.835 $X2=0.55 $Y2=2.91
r113 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.425
+ $Y=1.835 $X2=0.55 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%Y 1 2 3 4 5 6 7 8 27 33 35 36 37 38 41 47
+ 49 51 54 55 58 61 63 65 66 67 68 69 70 71 72 77 78
r148 78 80 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.2 $Y=0.97
+ $X2=4.44 $Y2=0.97
r149 77 86 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=5.39 $Y=0.97 $X2=5.3
+ $Y2=0.97
r150 72 77 4.35373 $w=4.3e-07 $l=1.3e-07 $layer=LI1_cond $X=5.52 $Y=0.97
+ $X2=5.39 $Y2=0.97
r151 71 86 6.96826 $w=4.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.04 $Y=0.97
+ $X2=5.3 $Y2=0.97
r152 70 71 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=0.97
+ $X2=5.04 $Y2=0.97
r153 70 80 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.56 $Y=0.97
+ $X2=4.44 $Y2=0.97
r154 69 78 4.58268 $w=4.3e-07 $l=1.40712e-07 $layer=LI1_cond $X=4.08 $Y=1.015
+ $X2=4.2 $Y2=0.97
r155 61 68 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=0.865
+ $X2=7.075 $Y2=0.865
r156 61 63 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=7.24 $Y=0.865
+ $X2=8.1 $Y2=0.865
r157 58 72 19.2488 $w=3.32e-07 $l=4.57329e-07 $layer=LI1_cond $X=5.965 $Y=0.945
+ $X2=5.52 $Y2=0.97
r158 58 68 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=5.965 $Y=0.945
+ $X2=7.075 $Y2=0.945
r159 56 67 5.0607 $w=2.05e-07 $l=3.51034e-07 $layer=LI1_cond $X=2.635 $Y=1.135
+ $X2=2.435 $Y2=0.87
r160 55 69 16.2998 $w=2.97e-07 $l=4.40936e-07 $layer=LI1_cond $X=3.695 $Y=1.135
+ $X2=4.08 $Y2=1.015
r161 55 56 50.8996 $w=2.38e-07 $l=1.06e-06 $layer=LI1_cond $X=3.695 $Y=1.135
+ $X2=2.635 $Y2=1.135
r162 53 67 1.43163 $w=2e-07 $l=4.32117e-07 $layer=LI1_cond $X=2.535 $Y=1.255
+ $X2=2.435 $Y2=0.87
r163 53 54 19.4091 $w=1.98e-07 $l=3.5e-07 $layer=LI1_cond $X=2.535 $Y=1.255
+ $X2=2.535 $Y2=1.605
r164 52 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.105 $Y=0.955
+ $X2=2.01 $Y2=0.955
r165 51 67 5.0607 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.955
+ $X2=2.435 $Y2=0.87
r166 51 52 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.435 $Y=0.955
+ $X2=2.105 $Y2=0.955
r167 50 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=1.69
+ $X2=1.84 $Y2=1.69
r168 49 54 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.435 $Y=1.69
+ $X2=2.535 $Y2=1.605
r169 49 50 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.435 $Y=1.69
+ $X2=2.005 $Y2=1.69
r170 45 66 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=0.87
+ $X2=2.01 $Y2=0.955
r171 45 47 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=2.01 $Y=0.87
+ $X2=2.01 $Y2=0.42
r172 41 43 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.84 $Y=1.96
+ $X2=1.84 $Y2=2.64
r173 39 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=1.775
+ $X2=1.84 $Y2=1.69
r174 39 41 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.84 $Y=1.775
+ $X2=1.84 $Y2=1.96
r175 37 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.915 $Y=0.955
+ $X2=2.01 $Y2=0.955
r176 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.915 $Y=0.955
+ $X2=1.245 $Y2=0.955
r177 35 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=1.69
+ $X2=1.84 $Y2=1.69
r178 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.675 $Y=1.69
+ $X2=1.145 $Y2=1.69
r179 31 38 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.15 $Y=0.87
+ $X2=1.245 $Y2=0.955
r180 31 33 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.15 $Y=0.87
+ $X2=1.15 $Y2=0.42
r181 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.98 $Y=1.96
+ $X2=0.98 $Y2=2.64
r182 25 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.98 $Y=1.775
+ $X2=1.145 $Y2=1.69
r183 25 27 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.98 $Y=1.775
+ $X2=0.98 $Y2=1.96
r184 8 43 400 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=1.7
+ $Y=1.835 $X2=1.84 $Y2=2.64
r185 8 41 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.7
+ $Y=1.835 $X2=1.84 $Y2=1.96
r186 7 29 400 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=0.84
+ $Y=1.835 $X2=0.98 $Y2=2.64
r187 7 27 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.84
+ $Y=1.835 $X2=0.98 $Y2=1.96
r188 6 63 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=7.96
+ $Y=0.235 $X2=8.1 $Y2=0.865
r189 5 61 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=7.1
+ $Y=0.235 $X2=7.24 $Y2=0.865
r190 4 86 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=5.16
+ $Y=0.235 $X2=5.3 $Y2=0.925
r191 3 80 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.235 $X2=4.44 $Y2=0.925
r192 2 47 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.235 $X2=2.01 $Y2=0.42
r193 1 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%A_533_367# 1 2 3 4 5 6 7 8 9 30 32 33 40 41
+ 47 48 49 52 54 58 60 63 66 68 69 72 80 82 84
c106 69 0 1.59281e-19 $X=9.055 $Y=1.69
c107 60 0 5.71875e-20 $X=8.795 $Y=2.04
r108 72 74 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=9.855 $Y=1.98
+ $X2=9.855 $Y2=2.91
r109 70 72 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=9.855 $Y=1.775
+ $X2=9.855 $Y2=1.98
r110 68 70 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.725 $Y=1.69
+ $X2=9.855 $Y2=1.775
r111 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.725 $Y=1.69
+ $X2=9.055 $Y2=1.69
r112 64 84 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=8.96 $Y=2.125
+ $X2=8.925 $Y2=2.04
r113 64 66 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=8.96 $Y=2.125
+ $X2=8.96 $Y2=2.44
r114 63 84 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.925 $Y=1.955
+ $X2=8.925 $Y2=2.04
r115 62 69 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=8.925 $Y=1.775
+ $X2=9.055 $Y2=1.69
r116 62 63 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=8.925 $Y=1.775
+ $X2=8.925 $Y2=1.955
r117 61 82 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.195 $Y=2.04
+ $X2=8.1 $Y2=2.04
r118 60 84 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.795 $Y=2.04
+ $X2=8.925 $Y2=2.04
r119 60 61 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.795 $Y=2.04
+ $X2=8.195 $Y2=2.04
r120 56 82 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.1 $Y=2.125
+ $X2=8.1 $Y2=2.04
r121 56 58 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=8.1 $Y=2.125
+ $X2=8.1 $Y2=2.475
r122 55 80 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.335 $Y=2.04
+ $X2=7.235 $Y2=2.04
r123 54 82 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.005 $Y=2.04
+ $X2=8.1 $Y2=2.04
r124 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.005 $Y=2.04
+ $X2=7.335 $Y2=2.04
r125 50 80 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=2.125
+ $X2=7.235 $Y2=2.04
r126 50 52 19.4091 $w=1.98e-07 $l=3.5e-07 $layer=LI1_cond $X=7.235 $Y=2.125
+ $X2=7.235 $Y2=2.475
r127 48 80 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.135 $Y=2.04
+ $X2=7.235 $Y2=2.04
r128 48 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.135 $Y=2.04
+ $X2=6.455 $Y2=2.04
r129 47 76 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=6.355 $Y=2.15
+ $X2=6.355 $Y2=2.27
r130 44 49 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.355 $Y=2.125
+ $X2=6.455 $Y2=2.04
r131 44 47 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=6.355 $Y=2.125
+ $X2=6.355 $Y2=2.15
r132 41 78 3.32334 $w=3.2e-07 $l=1.52e-07 $layer=LI1_cond $X=6.295 $Y=2.77
+ $X2=6.295 $Y2=2.922
r133 41 43 9.3636 $w=3.18e-07 $l=2.6e-07 $layer=LI1_cond $X=6.295 $Y=2.77
+ $X2=6.295 $Y2=2.51
r134 40 76 7.37399 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=6.295 $Y=2.43
+ $X2=6.295 $Y2=2.27
r135 40 43 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=6.295 $Y=2.43
+ $X2=6.295 $Y2=2.51
r136 37 39 32.4951 $w=3.03e-07 $l=8.6e-07 $layer=LI1_cond $X=4.51 $Y=2.922
+ $X2=5.37 $Y2=2.922
r137 35 37 32.4951 $w=3.03e-07 $l=8.6e-07 $layer=LI1_cond $X=3.65 $Y=2.922
+ $X2=4.51 $Y2=2.922
r138 33 35 26.2606 $w=3.03e-07 $l=6.95e-07 $layer=LI1_cond $X=2.955 $Y=2.922
+ $X2=3.65 $Y2=2.922
r139 32 78 3.49826 $w=3.05e-07 $l=1.6e-07 $layer=LI1_cond $X=6.135 $Y=2.922
+ $X2=6.295 $Y2=2.922
r140 32 39 28.9055 $w=3.03e-07 $l=7.65e-07 $layer=LI1_cond $X=6.135 $Y=2.922
+ $X2=5.37 $Y2=2.922
r141 28 33 6.83024 $w=3.05e-07 $l=2.28703e-07 $layer=LI1_cond $X=2.79 $Y=2.77
+ $X2=2.955 $Y2=2.922
r142 28 30 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.79 $Y=2.77
+ $X2=2.79 $Y2=2.39
r143 9 74 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=2.91
r144 9 72 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=1.98
r145 8 84 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.82
+ $Y=1.835 $X2=8.96 $Y2=1.98
r146 8 66 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=8.82
+ $Y=1.835 $X2=8.96 $Y2=2.44
r147 7 82 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.96
+ $Y=1.835 $X2=8.1 $Y2=2.04
r148 7 58 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=7.96
+ $Y=1.835 $X2=8.1 $Y2=2.475
r149 6 80 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=2.04
r150 6 52 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=2.475
r151 5 78 600 $w=1.7e-07 $l=1.17074e-06 $layer=licon1_PDIFF $count=1 $X=6.09
+ $Y=1.835 $X2=6.29 $Y2=2.91
r152 5 47 600 $w=1.7e-07 $l=4.25588e-07 $layer=licon1_PDIFF $count=1 $X=6.09
+ $Y=1.835 $X2=6.35 $Y2=2.15
r153 5 43 600 $w=1.7e-07 $l=7.68521e-07 $layer=licon1_PDIFF $count=1 $X=6.09
+ $Y=1.835 $X2=6.29 $Y2=2.51
r154 4 39 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.23
+ $Y=1.835 $X2=5.37 $Y2=2.91
r155 3 37 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.835 $X2=4.51 $Y2=2.91
r156 2 35 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.51
+ $Y=1.835 $X2=3.65 $Y2=2.91
r157 1 30 300 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.835 $X2=2.79 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%VPWR 1 2 3 4 15 19 21 25 29 34 35 36 37 38
+ 50 57 58 61 64
r119 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r120 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r121 58 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r122 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r123 55 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.555 $Y=3.33
+ $X2=9.39 $Y2=3.33
r124 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.555 $Y=3.33
+ $X2=9.84 $Y2=3.33
r125 54 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r126 54 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r127 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r128 51 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.53 $Y2=3.33
r129 51 53 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.88 $Y2=3.33
r130 50 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=9.39 $Y2=3.33
r131 50 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 49 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r133 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r134 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r135 45 46 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r136 41 45 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r137 41 42 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r138 38 46 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 38 42 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 36 48 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.505 $Y=3.33
+ $X2=7.44 $Y2=3.33
r141 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=3.33
+ $X2=7.67 $Y2=3.33
r142 34 45 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.48 $Y2=3.33
r143 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.79 $Y2=3.33
r144 33 48 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=7.44 $Y2=3.33
r145 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.79 $Y2=3.33
r146 29 32 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=9.39 $Y=2.03
+ $X2=9.39 $Y2=2.95
r147 27 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=3.33
r148 27 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=2.95
r149 23 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=3.245
+ $X2=8.53 $Y2=3.33
r150 23 25 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=8.53 $Y=3.245
+ $X2=8.53 $Y2=2.4
r151 22 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.67 $Y2=3.33
r152 21 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=8.53 $Y2=3.33
r153 21 22 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=7.835 $Y2=3.33
r154 17 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=3.33
r155 17 19 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=2.4
r156 13 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.79 $Y=3.245
+ $X2=6.79 $Y2=3.33
r157 13 15 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=6.79 $Y=3.245
+ $X2=6.79 $Y2=2.4
r158 4 32 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.25
+ $Y=1.835 $X2=9.39 $Y2=2.95
r159 4 29 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=9.25
+ $Y=1.835 $X2=9.39 $Y2=2.03
r160 3 25 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=8.39
+ $Y=1.835 $X2=8.53 $Y2=2.4
r161 2 19 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=7.53
+ $Y=1.835 $X2=7.67 $Y2=2.4
r162 1 15 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=6.64
+ $Y=1.835 $X2=6.79 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 51 52 54 55 57 58 60 61 62 64 85 92 98 101 105
r137 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r138 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r139 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r140 96 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r141 96 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r142 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r143 93 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=8.96 $Y2=0
r144 93 95 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=9.36 $Y2=0
r145 92 104 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=9.655 $Y=0
+ $X2=9.867 $Y2=0
r146 92 95 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.655 $Y=0 $X2=9.36
+ $Y2=0
r147 91 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r148 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r149 88 91 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r150 87 90 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r151 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r152 85 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.96 $Y2=0
r153 85 90 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.4
+ $Y2=0
r154 84 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r155 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r156 80 83 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6
+ $Y2=0
r157 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r158 78 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r159 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r160 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r161 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r162 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r163 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r164 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r165 69 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.72
+ $Y2=0
r166 69 71 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.2
+ $Y2=0
r167 67 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r168 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r169 64 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.72
+ $Y2=0
r170 64 66 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0
+ $X2=0.24 $Y2=0
r171 62 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r172 62 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r173 60 83 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.135 $Y=0 $X2=6
+ $Y2=0
r174 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.135 $Y=0 $X2=6.3
+ $Y2=0
r175 59 87 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.465 $Y=0 $X2=6.48
+ $Y2=0
r176 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.465 $Y=0 $X2=6.3
+ $Y2=0
r177 57 77 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.12
+ $Y2=0
r178 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.3
+ $Y2=0
r179 56 80 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.6
+ $Y2=0
r180 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.3
+ $Y2=0
r181 54 74 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.275 $Y=0
+ $X2=2.16 $Y2=0
r182 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.44
+ $Y2=0
r183 53 77 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.605 $Y=0
+ $X2=3.12 $Y2=0
r184 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=2.44
+ $Y2=0
r185 51 71 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.2
+ $Y2=0
r186 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.58
+ $Y2=0
r187 50 74 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.745 $Y=0
+ $X2=2.16 $Y2=0
r188 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.58
+ $Y2=0
r189 46 104 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=9.82 $Y=0.085
+ $X2=9.867 $Y2=0
r190 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.82 $Y=0.085
+ $X2=9.82 $Y2=0.38
r191 42 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0
r192 42 44 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0.575
r193 38 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=0.085 $X2=6.3
+ $Y2=0
r194 38 40 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.3 $Y=0.085
+ $X2=6.3 $Y2=0.565
r195 34 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.085 $X2=3.3
+ $Y2=0
r196 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0.38
r197 30 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.085
+ $X2=2.44 $Y2=0
r198 30 32 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.44 $Y=0.085
+ $X2=2.44 $Y2=0.575
r199 26 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r200 26 28 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.575
r201 22 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r202 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.38
r203 7 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.68
+ $Y=0.235 $X2=9.82 $Y2=0.38
r204 6 44 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=8.82
+ $Y=0.235 $X2=8.96 $Y2=0.575
r205 5 40 182 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_NDIFF $count=1 $X=6.16
+ $Y=0.235 $X2=6.3 $Y2=0.565
r206 4 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.16
+ $Y=0.235 $X2=3.3 $Y2=0.38
r207 3 32 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.235 $X2=2.44 $Y2=0.575
r208 2 28 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.58 $Y2=0.575
r209 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.72 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%A_546_47# 1 2 3 4 13 19 22 27
r36 27 29 20.9495 $w=1.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.725 $Y=0.42
+ $X2=3.725 $Y2=0.76
r37 22 24 5.25359 $w=1.88e-07 $l=9e-08 $layer=LI1_cond $X=2.87 $Y=0.67 $X2=2.87
+ $Y2=0.76
r38 17 19 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=4.87 $Y=0.42 $X2=5.87
+ $Y2=0.42
r39 17 27 36.8433 $w=3.28e-07 $l=1.055e-06 $layer=LI1_cond $X=4.87 $Y=0.42
+ $X2=3.815 $Y2=0.42
r40 14 24 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.965 $Y=0.76 $X2=2.87
+ $Y2=0.76
r41 13 29 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.635 $Y=0.76 $X2=3.725
+ $Y2=0.76
r42 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.635 $Y=0.76
+ $X2=2.965 $Y2=0.76
r43 4 19 182 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_NDIFF $count=1 $X=5.59
+ $Y=0.235 $X2=5.87 $Y2=0.42
r44 3 17 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.73
+ $Y=0.235 $X2=4.87 $Y2=0.42
r45 2 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.235 $X2=3.73 $Y2=0.42
r46 1 22 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.235 $X2=2.87 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_4%A_1334_47# 1 2 3 4 13 19 20 21 25
c30 13 0 1.1786e-19 $X=8.425 $Y=0.392
r31 23 25 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=9.39 $Y=0.87
+ $X2=9.39 $Y2=0.42
r32 22 30 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.625 $Y=0.955
+ $X2=8.525 $Y2=0.955
r33 21 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=9.295 $Y=0.955
+ $X2=9.39 $Y2=0.87
r34 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.295 $Y=0.955
+ $X2=8.625 $Y2=0.955
r35 20 30 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=0.87 $X2=8.525
+ $Y2=0.955
r36 19 28 4.08194 $w=2e-07 $l=1.38e-07 $layer=LI1_cond $X=8.525 $Y=0.53
+ $X2=8.525 $Y2=0.392
r37 19 20 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=8.525 $Y=0.53
+ $X2=8.525 $Y2=0.87
r38 15 18 36.04 $w=2.73e-07 $l=8.6e-07 $layer=LI1_cond $X=6.81 $Y=0.392 $X2=7.67
+ $Y2=0.392
r39 13 28 2.95793 $w=2.75e-07 $l=1e-07 $layer=LI1_cond $X=8.425 $Y=0.392
+ $X2=8.525 $Y2=0.392
r40 13 18 31.6398 $w=2.73e-07 $l=7.55e-07 $layer=LI1_cond $X=8.425 $Y=0.392
+ $X2=7.67 $Y2=0.392
r41 4 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.25
+ $Y=0.235 $X2=9.39 $Y2=0.42
r42 3 30 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=8.39
+ $Y=0.235 $X2=8.53 $Y2=0.875
r43 3 28 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=8.39
+ $Y=0.235 $X2=8.53 $Y2=0.42
r44 2 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.53
+ $Y=0.235 $X2=7.67 $Y2=0.38
r45 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.67
+ $Y=0.235 $X2=6.81 $Y2=0.38
.ends

