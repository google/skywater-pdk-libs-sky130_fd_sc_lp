* NGSPICE file created from sky130_fd_sc_lp__iso0n_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__iso0n_lp2 A SLEEP_B KAGND VGND VNB VPB VPWR X
M1000 VPWR SLEEP_B a_65_65# VPB phighvt w=1e+06u l=250000u
+  ad=6.3e+11p pd=5.26e+06u as=2.8e+11p ps=2.56e+06u
M1001 a_152_65# A a_65_65# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1002 KAGND SLEEP_B a_152_65# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1003 X a_65_65# a_316_65# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_316_65# a_65_65# KAGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_65_65# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_65_65# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

