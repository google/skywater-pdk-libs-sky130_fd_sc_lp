* File: sky130_fd_sc_lp__fa_0.pxi.spice
* Created: Fri Aug 28 10:34:35 2020
* 
x_PM_SKY130_FD_SC_LP__FA_0%A N_A_M1010_g N_A_M1003_g N_A_c_162_n N_A_c_163_n
+ N_A_M1016_g N_A_M1023_g N_A_c_164_n N_A_c_165_n N_A_c_166_n N_A_c_167_n
+ N_A_M1013_g N_A_M1008_g N_A_c_169_n N_A_M1001_g N_A_M1015_g N_A_c_171_n
+ N_A_c_172_n N_A_c_156_n N_A_c_157_n N_A_c_174_n A A A N_A_c_158_n N_A_c_159_n
+ PM_SKY130_FD_SC_LP__FA_0%A
x_PM_SKY130_FD_SC_LP__FA_0%B N_B_M1020_g N_B_M1025_g N_B_M1027_g N_B_M1021_g
+ N_B_M1017_g N_B_M1018_g N_B_M1014_g N_B_c_328_n N_B_M1009_g N_B_c_329_n
+ N_B_c_330_n N_B_c_340_n N_B_c_341_n N_B_c_342_n N_B_c_343_n N_B_c_344_n
+ N_B_c_345_n B B B N_B_c_332_n PM_SKY130_FD_SC_LP__FA_0%B
x_PM_SKY130_FD_SC_LP__FA_0%CIN N_CIN_M1022_g N_CIN_M1005_g N_CIN_M1002_g
+ N_CIN_M1004_g N_CIN_M1012_g N_CIN_M1019_g N_CIN_c_496_n N_CIN_c_497_n
+ N_CIN_c_498_n N_CIN_c_499_n N_CIN_c_500_n CIN N_CIN_c_501_n N_CIN_c_502_n
+ PM_SKY130_FD_SC_LP__FA_0%CIN
x_PM_SKY130_FD_SC_LP__FA_0%A_80_225# N_A_80_225#_M1020_d N_A_80_225#_M1025_d
+ N_A_80_225#_M1007_g N_A_80_225#_M1026_g N_A_80_225#_c_612_n
+ N_A_80_225#_c_613_n N_A_80_225#_M1011_g N_A_80_225#_M1024_g
+ N_A_80_225#_c_616_n N_A_80_225#_c_617_n N_A_80_225#_c_618_n
+ N_A_80_225#_c_625_n N_A_80_225#_c_626_n N_A_80_225#_c_627_n
+ N_A_80_225#_c_653_n N_A_80_225#_c_667_n N_A_80_225#_c_619_n
+ N_A_80_225#_c_620_n N_A_80_225#_c_621_n N_A_80_225#_c_657_n
+ PM_SKY130_FD_SC_LP__FA_0%A_80_225#
x_PM_SKY130_FD_SC_LP__FA_0%A_1059_119# N_A_1059_119#_M1011_d
+ N_A_1059_119#_M1024_d N_A_1059_119#_M1006_g N_A_1059_119#_M1000_g
+ N_A_1059_119#_c_741_n N_A_1059_119#_c_754_n N_A_1059_119#_c_742_n
+ N_A_1059_119#_c_743_n N_A_1059_119#_c_759_n N_A_1059_119#_c_744_n
+ N_A_1059_119#_c_745_n N_A_1059_119#_c_746_n N_A_1059_119#_c_747_n
+ N_A_1059_119#_c_748_n PM_SKY130_FD_SC_LP__FA_0%A_1059_119#
x_PM_SKY130_FD_SC_LP__FA_0%COUT N_COUT_M1026_s N_COUT_M1007_s N_COUT_c_814_n
+ N_COUT_c_816_n COUT COUT COUT COUT PM_SKY130_FD_SC_LP__FA_0%COUT
x_PM_SKY130_FD_SC_LP__FA_0%VPWR N_VPWR_M1007_d N_VPWR_M1021_d N_VPWR_M1004_s
+ N_VPWR_M1018_d N_VPWR_M1015_d N_VPWR_c_832_n N_VPWR_c_833_n N_VPWR_c_834_n
+ N_VPWR_c_835_n N_VPWR_c_836_n VPWR N_VPWR_c_837_n N_VPWR_c_838_n
+ N_VPWR_c_839_n N_VPWR_c_840_n N_VPWR_c_841_n N_VPWR_c_842_n N_VPWR_c_831_n
+ N_VPWR_c_844_n N_VPWR_c_845_n N_VPWR_c_846_n N_VPWR_c_847_n N_VPWR_c_848_n
+ PM_SKY130_FD_SC_LP__FA_0%VPWR
x_PM_SKY130_FD_SC_LP__FA_0%A_404_532# N_A_404_532#_M1005_d N_A_404_532#_M1016_d
+ N_A_404_532#_c_936_n N_A_404_532#_c_928_n N_A_404_532#_c_929_n
+ N_A_404_532#_c_930_n PM_SKY130_FD_SC_LP__FA_0%A_404_532#
x_PM_SKY130_FD_SC_LP__FA_0%A_781_457# N_A_781_457#_M1004_d N_A_781_457#_M1008_d
+ N_A_781_457#_c_956_n N_A_781_457#_c_957_n N_A_781_457#_c_958_n
+ N_A_781_457#_c_959_n PM_SKY130_FD_SC_LP__FA_0%A_781_457#
x_PM_SKY130_FD_SC_LP__FA_0%SUM N_SUM_M1006_d N_SUM_M1000_d N_SUM_c_987_n
+ N_SUM_c_988_n SUM SUM SUM SUM SUM SUM PM_SKY130_FD_SC_LP__FA_0%SUM
x_PM_SKY130_FD_SC_LP__FA_0%VGND N_VGND_M1026_d N_VGND_M1027_d N_VGND_M1002_s
+ N_VGND_M1017_d N_VGND_M1001_d N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n VGND
+ N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n
+ N_VGND_c_1015_n N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n
+ N_VGND_c_1019_n PM_SKY130_FD_SC_LP__FA_0%VGND
x_PM_SKY130_FD_SC_LP__FA_0%A_382_119# N_A_382_119#_M1022_d N_A_382_119#_M1023_d
+ N_A_382_119#_c_1096_n N_A_382_119#_c_1097_n N_A_382_119#_c_1098_n
+ PM_SKY130_FD_SC_LP__FA_0%A_382_119#
x_PM_SKY130_FD_SC_LP__FA_0%A_781_119# N_A_781_119#_M1002_d N_A_781_119#_M1013_d
+ N_A_781_119#_c_1125_n N_A_781_119#_c_1123_n N_A_781_119#_c_1124_n
+ N_A_781_119#_c_1127_n PM_SKY130_FD_SC_LP__FA_0%A_781_119#
cc_1 VNB N_A_M1003_g 0.0381415f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.805
cc_2 VNB N_A_M1023_g 0.0421138f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.805
cc_3 VNB N_A_M1013_g 0.0420894f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=0.805
cc_4 VNB N_A_M1001_g 0.0494439f $X=-0.19 $Y=-0.245 $X2=6.64 $Y2=0.515
cc_5 VNB N_A_M1015_g 0.00596245f $X=-0.19 $Y=-0.245 $X2=6.66 $Y2=2.495
cc_6 VNB N_A_c_156_n 0.0114921f $X=-0.19 $Y=-0.245 $X2=6.665 $Y2=1.555
cc_7 VNB N_A_c_157_n 0.00166459f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.695
cc_8 VNB N_A_c_158_n 0.0160954f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=1.665
cc_9 VNB N_A_c_159_n 0.0137623f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=1.665
cc_10 VNB N_B_M1020_g 0.0374407f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.87
cc_11 VNB N_B_M1017_g 0.0423749f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=2.55
cc_12 VNB N_B_M1014_g 0.0420102f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=2.495
cc_13 VNB N_B_c_328_n 0.00452492f $X=-0.19 $Y=-0.245 $X2=6.585 $Y2=3.15
cc_14 VNB N_B_c_329_n 0.0162414f $X=-0.19 $Y=-0.245 $X2=6.64 $Y2=0.515
cc_15 VNB N_B_c_330_n 0.00989428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB B 0.00413984f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_17 VNB N_B_c_332_n 0.0177981f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=1.5
cc_18 VNB N_CIN_M1022_g 0.0171998f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.87
cc_19 VNB N_CIN_M1005_g 0.00886044f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.805
cc_20 VNB N_CIN_M1002_g 0.0242124f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.55
cc_21 VNB N_CIN_M1004_g 0.00830645f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.805
cc_22 VNB N_CIN_M1012_g 0.0271354f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=2.475
cc_23 VNB N_CIN_M1019_g 0.00160942f $X=-0.19 $Y=-0.245 $X2=3.415 $Y2=3.15
cc_24 VNB N_CIN_c_496_n 0.0290172f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=0.805
cc_25 VNB N_CIN_c_497_n 0.0301241f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=2.495
cc_26 VNB N_CIN_c_498_n 0.00289181f $X=-0.19 $Y=-0.245 $X2=6.64 $Y2=0.515
cc_27 VNB N_CIN_c_499_n 0.0280119f $X=-0.19 $Y=-0.245 $X2=6.64 $Y2=0.515
cc_28 VNB N_CIN_c_500_n 0.0230975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_CIN_c_501_n 0.00969258f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.695
cc_30 VNB N_CIN_c_502_n 0.0472947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_80_225#_M1007_g 0.0110216f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.83
cc_32 VNB N_A_80_225#_M1026_g 0.0353855f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=1.5
cc_33 VNB N_A_80_225#_c_612_n 0.339915f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.805
cc_34 VNB N_A_80_225#_c_613_n 0.0126405f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.805
cc_35 VNB N_A_80_225#_M1011_g 0.0317071f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=2.55
cc_36 VNB N_A_80_225#_M1024_g 0.0170731f $X=-0.19 $Y=-0.245 $X2=3.415 $Y2=3.15
cc_37 VNB N_A_80_225#_c_616_n 0.00961548f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=0.805
cc_38 VNB N_A_80_225#_c_617_n 0.00171482f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=2.495
cc_39 VNB N_A_80_225#_c_618_n 0.0137883f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=2.495
cc_40 VNB N_A_80_225#_c_619_n 0.0021364f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.475
cc_41 VNB N_A_80_225#_c_620_n 0.00175969f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=3.15
cc_42 VNB N_A_80_225#_c_621_n 0.0370856f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.695
cc_43 VNB N_A_1059_119#_M1000_g 0.0274711f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.87
cc_44 VNB N_A_1059_119#_c_741_n 0.0101855f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=1.5
cc_45 VNB N_A_1059_119#_c_742_n 0.00603143f $X=-0.19 $Y=-0.245 $X2=3.34
+ $Y2=3.075
cc_46 VNB N_A_1059_119#_c_743_n 0.00293298f $X=-0.19 $Y=-0.245 $X2=3.415
+ $Y2=3.15
cc_47 VNB N_A_1059_119#_c_744_n 0.00212215f $X=-0.19 $Y=-0.245 $X2=6.64
+ $Y2=1.405
cc_48 VNB N_A_1059_119#_c_745_n 0.00175621f $X=-0.19 $Y=-0.245 $X2=6.64
+ $Y2=0.515
cc_49 VNB N_A_1059_119#_c_746_n 0.00380798f $X=-0.19 $Y=-0.245 $X2=6.66
+ $Y2=1.555
cc_50 VNB N_A_1059_119#_c_747_n 0.0416007f $X=-0.19 $Y=-0.245 $X2=6.66 $Y2=3.075
cc_51 VNB N_A_1059_119#_c_748_n 0.0207586f $X=-0.19 $Y=-0.245 $X2=2.845
+ $Y2=2.475
cc_52 VNB N_COUT_c_814_n 0.0178523f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.87
cc_53 VNB COUT 0.0357991f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=2.475
cc_54 VNB N_VPWR_c_831_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SUM_c_987_n 0.0170074f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.4
cc_56 VNB N_SUM_c_988_n 0.00953258f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=1.5
cc_57 VNB SUM 0.0377987f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.805
cc_58 VNB SUM 0.00566811f $X=-0.19 $Y=-0.245 $X2=3.265 $Y2=2.475
cc_59 VNB N_VGND_c_1004_n 0.00831555f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=2.55
cc_60 VNB N_VGND_c_1005_n 0.0191927f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=3.075
cc_61 VNB N_VGND_c_1006_n 0.0176618f $X=-0.19 $Y=-0.245 $X2=4.79 $Y2=2.495
cc_62 VNB N_VGND_c_1007_n 0.0102682f $X=-0.19 $Y=-0.245 $X2=6.64 $Y2=1.405
cc_63 VNB N_VGND_c_1008_n 0.00447809f $X=-0.19 $Y=-0.245 $X2=6.66 $Y2=1.555
cc_64 VNB N_VGND_c_1009_n 0.0593695f $X=-0.19 $Y=-0.245 $X2=6.66 $Y2=2.495
cc_65 VNB N_VGND_c_1010_n 0.00499185f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.475
cc_66 VNB N_VGND_c_1011_n 0.0394288f $X=-0.19 $Y=-0.245 $X2=6.665 $Y2=1.555
cc_67 VNB N_VGND_c_1012_n 0.0188756f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_68 VNB N_VGND_c_1013_n 0.0152411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1014_n 0.0208241f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.695
cc_70 VNB N_VGND_c_1015_n 0.39397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1016_n 0.0247945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1017_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1018_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1019_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_382_119#_c_1096_n 0.00327133f $X=-0.19 $Y=-0.245 $X2=1.045
+ $Y2=0.805
cc_76 VNB N_A_382_119#_c_1097_n 0.00309147f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.4
cc_77 VNB N_A_382_119#_c_1098_n 0.00782281f $X=-0.19 $Y=-0.245 $X2=2.855
+ $Y2=0.805
cc_78 VNB N_A_781_119#_c_1123_n 0.0115252f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=2.55
cc_79 VNB N_A_781_119#_c_1124_n 0.00373405f $X=-0.19 $Y=-0.245 $X2=2.845
+ $Y2=2.87
cc_80 VPB N_A_M1010_g 0.0430944f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.87
cc_81 VPB N_A_M1003_g 0.0017274f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.805
cc_82 VPB N_A_c_162_n 0.0332068f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.4
cc_83 VPB N_A_c_163_n 0.0160727f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.55
cc_84 VPB N_A_c_164_n 0.0284515f $X=-0.19 $Y=1.655 $X2=3.265 $Y2=2.475
cc_85 VPB N_A_c_165_n 0.0295798f $X=-0.19 $Y=1.655 $X2=3.34 $Y2=3.075
cc_86 VPB N_A_c_166_n 0.0903528f $X=-0.19 $Y=1.655 $X2=4.715 $Y2=3.15
cc_87 VPB N_A_c_167_n 0.0101954f $X=-0.19 $Y=1.655 $X2=3.415 $Y2=3.15
cc_88 VPB N_A_M1013_g 0.0581877f $X=-0.19 $Y=1.655 $X2=4.79 $Y2=0.805
cc_89 VPB N_A_c_169_n 0.137216f $X=-0.19 $Y=1.655 $X2=6.585 $Y2=3.15
cc_90 VPB N_A_M1015_g 0.064708f $X=-0.19 $Y=1.655 $X2=6.66 $Y2=2.495
cc_91 VPB N_A_c_171_n 0.00522616f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.475
cc_92 VPB N_A_c_172_n 0.00749069f $X=-0.19 $Y=1.655 $X2=4.79 $Y2=3.15
cc_93 VPB N_A_c_157_n 0.0011753f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.695
cc_94 VPB N_A_c_174_n 0.03201f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=1.86
cc_95 VPB N_A_c_158_n 0.0173014f $X=-0.19 $Y=1.655 $X2=2.785 $Y2=1.665
cc_96 VPB N_A_c_159_n 0.0165096f $X=-0.19 $Y=1.655 $X2=2.785 $Y2=1.665
cc_97 VPB N_B_M1020_g 0.01651f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.87
cc_98 VPB N_B_M1025_g 0.0302113f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.805
cc_99 VPB N_B_M1021_g 0.02321f $X=-0.19 $Y=1.655 $X2=2.855 $Y2=0.805
cc_100 VPB N_B_M1017_g 0.00109903f $X=-0.19 $Y=1.655 $X2=3.34 $Y2=2.55
cc_101 VPB N_B_M1018_g 0.0241903f $X=-0.19 $Y=1.655 $X2=4.79 $Y2=3.075
cc_102 VPB N_B_c_328_n 0.0353409f $X=-0.19 $Y=1.655 $X2=6.585 $Y2=3.15
cc_103 VPB N_B_M1009_g 0.019092f $X=-0.19 $Y=1.655 $X2=6.64 $Y2=1.405
cc_104 VPB N_B_c_340_n 0.0198209f $X=-0.19 $Y=1.655 $X2=6.66 $Y2=1.555
cc_105 VPB N_B_c_341_n 0.0301657f $X=-0.19 $Y=1.655 $X2=6.66 $Y2=2.495
cc_106 VPB N_B_c_342_n 0.0287311f $X=-0.19 $Y=1.655 $X2=6.665 $Y2=1.555
cc_107 VPB N_B_c_343_n 0.0541851f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.695
cc_108 VPB N_B_c_344_n 0.0296685f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=1.86
cc_109 VPB N_B_c_345_n 0.01468f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=1.86
cc_110 VPB B 5.93334e-19 $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.58
cc_111 VPB N_B_c_332_n 0.0190934f $X=-0.19 $Y=1.655 $X2=2.785 $Y2=1.5
cc_112 VPB N_CIN_M1005_g 0.0589953f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=0.805
cc_113 VPB N_CIN_M1004_g 0.049969f $X=-0.19 $Y=1.655 $X2=2.855 $Y2=0.805
cc_114 VPB N_CIN_M1019_g 0.0429561f $X=-0.19 $Y=1.655 $X2=3.415 $Y2=3.15
cc_115 VPB N_A_80_225#_M1007_g 0.055396f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=1.83
cc_116 VPB N_A_80_225#_M1024_g 0.0432327f $X=-0.19 $Y=1.655 $X2=3.415 $Y2=3.15
cc_117 VPB N_A_80_225#_c_617_n 0.00388859f $X=-0.19 $Y=1.655 $X2=4.79 $Y2=2.495
cc_118 VPB N_A_80_225#_c_625_n 0.0111542f $X=-0.19 $Y=1.655 $X2=4.865 $Y2=3.15
cc_119 VPB N_A_80_225#_c_626_n 0.00306875f $X=-0.19 $Y=1.655 $X2=6.64 $Y2=1.405
cc_120 VPB N_A_80_225#_c_627_n 0.00271241f $X=-0.19 $Y=1.655 $X2=6.64 $Y2=0.515
cc_121 VPB N_A_1059_119#_M1000_g 0.0514444f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.87
cc_122 VPB N_A_1059_119#_c_742_n 0.0122712f $X=-0.19 $Y=1.655 $X2=3.34 $Y2=3.075
cc_123 VPB N_COUT_c_816_n 0.0228675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB COUT 0.0419089f $X=-0.19 $Y=1.655 $X2=2.92 $Y2=2.475
cc_125 VPB N_VPWR_c_832_n 0.00641629f $X=-0.19 $Y=1.655 $X2=3.265 $Y2=2.475
cc_126 VPB N_VPWR_c_833_n 8.75318e-19 $X=-0.19 $Y=1.655 $X2=4.715 $Y2=3.15
cc_127 VPB N_VPWR_c_834_n 0.0132508f $X=-0.19 $Y=1.655 $X2=4.79 $Y2=0.805
cc_128 VPB N_VPWR_c_835_n 0.0107618f $X=-0.19 $Y=1.655 $X2=6.585 $Y2=3.15
cc_129 VPB N_VPWR_c_836_n 0.0110491f $X=-0.19 $Y=1.655 $X2=6.64 $Y2=0.515
cc_130 VPB N_VPWR_c_837_n 0.0177734f $X=-0.19 $Y=1.655 $X2=6.66 $Y2=2.495
cc_131 VPB N_VPWR_c_838_n 0.0386942f $X=-0.19 $Y=1.655 $X2=6.665 $Y2=1.555
cc_132 VPB N_VPWR_c_839_n 0.016926f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_133 VPB N_VPWR_c_840_n 0.016234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_841_n 0.0636179f $X=-0.19 $Y=1.655 $X2=2.785 $Y2=1.665
cc_135 VPB N_VPWR_c_842_n 0.0173857f $X=-0.19 $Y=1.655 $X2=2.785 $Y2=1.695
cc_136 VPB N_VPWR_c_831_n 0.069023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_844_n 0.00564503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_845_n 0.0045467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_846_n 0.00363625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_847_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_848_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_404_532#_c_928_n 0.00652549f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.55
cc_143 VPB N_A_404_532#_c_929_n 0.00222594f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.87
cc_144 VPB N_A_404_532#_c_930_n 0.00319287f $X=-0.19 $Y=1.655 $X2=2.855
+ $Y2=0.805
cc_145 VPB N_A_781_457#_c_956_n 2.27481e-19 $X=-0.19 $Y=1.655 $X2=2.845 $Y2=1.83
cc_146 VPB N_A_781_457#_c_957_n 0.0111411f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.55
cc_147 VPB N_A_781_457#_c_958_n 0.00452375f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=2.87
cc_148 VPB N_A_781_457#_c_959_n 2.40439e-19 $X=-0.19 $Y=1.655 $X2=2.855
+ $Y2=0.805
cc_149 VPB SUM 0.0628163f $X=-0.19 $Y=1.655 $X2=3.265 $Y2=2.475
cc_150 N_A_M1003_g N_B_M1020_g 0.0482608f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_151 N_A_c_157_n N_B_M1020_g 0.00143509f $X=0.995 $Y=1.695 $X2=0 $Y2=0
cc_152 N_A_c_159_n N_B_M1020_g 0.0165052f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_153 N_A_c_171_n N_B_M1021_g 0.0185652f $X=2.845 $Y=2.475 $X2=0 $Y2=0
cc_154 N_A_M1013_g N_B_M1017_g 0.0271116f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_155 N_A_c_166_n N_B_M1018_g 0.00907339f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_156 N_A_M1013_g N_B_M1018_g 0.0136931f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_157 N_A_M1001_g N_B_M1014_g 0.0364045f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_158 N_A_M1015_g N_B_M1014_g 7.24147e-19 $X=6.66 $Y=2.495 $X2=0 $Y2=0
cc_159 N_A_M1015_g N_B_c_328_n 0.0251681f $X=6.66 $Y=2.495 $X2=0 $Y2=0
cc_160 N_A_c_169_n N_B_M1009_g 0.00865213f $X=6.585 $Y=3.15 $X2=0 $Y2=0
cc_161 N_A_M1015_g N_B_M1009_g 0.0234897f $X=6.66 $Y=2.495 $X2=0 $Y2=0
cc_162 N_A_M1023_g N_B_c_329_n 0.0168299f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_163 N_A_M1023_g N_B_c_330_n 0.0134073f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_164 N_A_M1010_g N_B_c_340_n 0.00104017f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_165 N_A_c_162_n N_B_c_340_n 0.0182493f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_c_164_n N_B_c_340_n 0.00477753f $X=3.265 $Y=2.475 $X2=0 $Y2=0
cc_167 N_A_c_157_n N_B_c_340_n 0.00178228f $X=0.995 $Y=1.695 $X2=0 $Y2=0
cc_168 N_A_c_158_n N_B_c_340_n 0.00377412f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_169 N_A_c_159_n N_B_c_340_n 0.120671f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_170 N_A_M1010_g N_B_c_341_n 0.0626465f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_171 N_A_c_174_n N_B_c_341_n 0.0482608f $X=0.955 $Y=1.86 $X2=0 $Y2=0
cc_172 N_A_c_159_n N_B_c_341_n 0.00407239f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_173 N_A_c_162_n N_B_c_342_n 0.0217391f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_c_159_n N_B_c_342_n 0.00105694f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_175 N_A_c_164_n N_B_c_343_n 0.00346402f $X=3.265 $Y=2.475 $X2=0 $Y2=0
cc_176 N_A_M1013_g N_B_c_343_n 0.0101493f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_177 N_A_M1013_g N_B_c_344_n 0.0192649f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_178 N_A_c_162_n N_B_c_345_n 0.00670205f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_c_164_n N_B_c_345_n 0.00629517f $X=3.265 $Y=2.475 $X2=0 $Y2=0
cc_180 N_A_c_158_n N_B_c_345_n 8.54377e-19 $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_181 N_A_c_159_n N_B_c_345_n 0.00489697f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_182 N_A_M1001_g B 0.00540955f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_183 N_A_M1015_g B 0.00481823f $X=6.66 $Y=2.495 $X2=0 $Y2=0
cc_184 N_A_c_156_n B 0.00457874f $X=6.665 $Y=1.555 $X2=0 $Y2=0
cc_185 N_A_c_162_n N_B_c_332_n 0.00902743f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A_c_158_n N_B_c_332_n 0.0217775f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_187 N_A_c_159_n N_B_c_332_n 0.0124249f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_188 N_A_c_159_n N_CIN_M1005_g 0.0139333f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_189 N_A_c_164_n N_CIN_M1004_g 0.00815451f $X=3.265 $Y=2.475 $X2=0 $Y2=0
cc_190 N_A_c_166_n N_CIN_M1004_g 0.00907339f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_191 N_A_c_169_n N_CIN_M1019_g 0.00865213f $X=6.585 $Y=3.15 $X2=0 $Y2=0
cc_192 N_A_M1023_g N_CIN_c_496_n 0.0118687f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_193 N_A_c_158_n N_CIN_c_496_n 0.00442627f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_194 N_A_c_159_n N_CIN_c_496_n 0.0928664f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_195 N_A_c_159_n N_CIN_c_497_n 0.00495247f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_196 N_A_M1013_g N_CIN_c_500_n 0.0129954f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_197 N_A_M1023_g N_CIN_c_501_n 0.00269997f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_198 N_A_c_158_n N_CIN_c_501_n 0.00132325f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_199 N_A_c_159_n N_CIN_c_501_n 5.6664e-19 $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_200 N_A_M1023_g N_CIN_c_502_n 0.0056572f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_201 N_A_c_158_n N_CIN_c_502_n 8.50415e-19 $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_202 N_A_M1010_g N_A_80_225#_M1007_g 0.0227226f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_203 N_A_M1003_g N_A_80_225#_M1007_g 0.00586761f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_204 N_A_c_157_n N_A_80_225#_M1007_g 6.13597e-19 $X=0.995 $Y=1.695 $X2=0 $Y2=0
cc_205 N_A_c_174_n N_A_80_225#_M1007_g 0.0171216f $X=0.955 $Y=1.86 $X2=0 $Y2=0
cc_206 N_A_M1003_g N_A_80_225#_M1026_g 0.0119911f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_207 N_A_M1003_g N_A_80_225#_c_612_n 0.0103107f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_208 N_A_M1023_g N_A_80_225#_c_612_n 0.0100733f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_209 N_A_M1013_g N_A_80_225#_c_612_n 0.0104164f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_210 N_A_M1013_g N_A_80_225#_M1011_g 0.0115947f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_211 N_A_M1013_g N_A_80_225#_M1024_g 0.0548831f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_212 N_A_c_169_n N_A_80_225#_M1024_g 0.00907339f $X=6.585 $Y=3.15 $X2=0 $Y2=0
cc_213 N_A_M1013_g N_A_80_225#_c_616_n 0.00820047f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_214 N_A_M1010_g N_A_80_225#_c_617_n 0.00337916f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_215 N_A_M1003_g N_A_80_225#_c_617_n 0.00257517f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_216 N_A_c_157_n N_A_80_225#_c_617_n 0.0339783f $X=0.995 $Y=1.695 $X2=0 $Y2=0
cc_217 N_A_c_174_n N_A_80_225#_c_617_n 0.00220024f $X=0.955 $Y=1.86 $X2=0 $Y2=0
cc_218 N_A_M1003_g N_A_80_225#_c_618_n 0.0137789f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_219 N_A_c_157_n N_A_80_225#_c_618_n 0.0132435f $X=0.995 $Y=1.695 $X2=0 $Y2=0
cc_220 N_A_c_174_n N_A_80_225#_c_618_n 0.00287367f $X=0.955 $Y=1.86 $X2=0 $Y2=0
cc_221 N_A_c_159_n N_A_80_225#_c_618_n 0.021726f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_222 N_A_M1010_g N_A_80_225#_c_625_n 0.0132639f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_223 N_A_c_157_n N_A_80_225#_c_625_n 0.0191259f $X=0.995 $Y=1.695 $X2=0 $Y2=0
cc_224 N_A_c_174_n N_A_80_225#_c_625_n 0.00375607f $X=0.955 $Y=1.86 $X2=0 $Y2=0
cc_225 N_A_c_159_n N_A_80_225#_c_625_n 0.0055104f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_226 N_A_M1010_g N_A_80_225#_c_627_n 0.00832821f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_227 N_A_M1010_g N_A_80_225#_c_653_n 0.00720972f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_228 N_A_M1003_g N_A_80_225#_c_619_n 0.00349968f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_229 N_A_M1003_g N_A_80_225#_c_620_n 0.0010329f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_230 N_A_M1003_g N_A_80_225#_c_621_n 0.0208532f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_231 N_A_M1003_g N_A_80_225#_c_657_n 0.00261393f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_232 N_A_c_159_n N_A_80_225#_c_657_n 0.00523018f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_233 N_A_M1001_g N_A_1059_119#_M1000_g 0.00413049f $X=6.64 $Y=0.515 $X2=0
+ $Y2=0
cc_234 N_A_M1015_g N_A_1059_119#_M1000_g 0.0301905f $X=6.66 $Y=2.495 $X2=0 $Y2=0
cc_235 N_A_c_156_n N_A_1059_119#_M1000_g 0.00422554f $X=6.665 $Y=1.555 $X2=0
+ $Y2=0
cc_236 N_A_c_169_n N_A_1059_119#_c_754_n 0.0108101f $X=6.585 $Y=3.15 $X2=0 $Y2=0
cc_237 N_A_M1015_g N_A_1059_119#_c_754_n 0.0200786f $X=6.66 $Y=2.495 $X2=0 $Y2=0
cc_238 N_A_M1001_g N_A_1059_119#_c_742_n 0.00194193f $X=6.64 $Y=0.515 $X2=0
+ $Y2=0
cc_239 N_A_M1015_g N_A_1059_119#_c_742_n 0.00986295f $X=6.66 $Y=2.495 $X2=0
+ $Y2=0
cc_240 N_A_c_156_n N_A_1059_119#_c_742_n 0.00459241f $X=6.665 $Y=1.555 $X2=0
+ $Y2=0
cc_241 N_A_c_169_n N_A_1059_119#_c_759_n 0.00553204f $X=6.585 $Y=3.15 $X2=0
+ $Y2=0
cc_242 N_A_M1001_g N_A_1059_119#_c_744_n 4.64877e-19 $X=6.64 $Y=0.515 $X2=0
+ $Y2=0
cc_243 N_A_M1001_g N_A_1059_119#_c_745_n 0.0159408f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_244 N_A_c_156_n N_A_1059_119#_c_745_n 9.19703e-19 $X=6.665 $Y=1.555 $X2=0
+ $Y2=0
cc_245 N_A_M1001_g N_A_1059_119#_c_746_n 0.00495926f $X=6.64 $Y=0.515 $X2=0
+ $Y2=0
cc_246 N_A_M1001_g N_A_1059_119#_c_747_n 0.0221857f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_247 N_A_M1001_g N_A_1059_119#_c_748_n 0.0122468f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_248 N_A_M1010_g N_COUT_c_816_n 5.85497e-19 $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_249 N_A_M1010_g N_VPWR_c_832_n 0.00332345f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_250 N_A_c_163_n N_VPWR_c_833_n 0.00687623f $X=2.845 $Y=2.55 $X2=0 $Y2=0
cc_251 N_A_c_165_n N_VPWR_c_833_n 0.00117131f $X=3.34 $Y=3.075 $X2=0 $Y2=0
cc_252 N_A_c_167_n N_VPWR_c_833_n 2.65719e-19 $X=3.415 $Y=3.15 $X2=0 $Y2=0
cc_253 N_A_c_162_n N_VPWR_c_834_n 0.0018184f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A_c_163_n N_VPWR_c_834_n 7.90819e-19 $X=2.845 $Y=2.55 $X2=0 $Y2=0
cc_255 N_A_c_164_n N_VPWR_c_834_n 0.0122399f $X=3.265 $Y=2.475 $X2=0 $Y2=0
cc_256 N_A_c_166_n N_VPWR_c_834_n 0.0206256f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_257 N_A_c_166_n N_VPWR_c_835_n 0.0236268f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_258 N_A_M1013_g N_VPWR_c_835_n 0.0142225f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_259 N_A_M1015_g N_VPWR_c_836_n 0.0182662f $X=6.66 $Y=2.495 $X2=0 $Y2=0
cc_260 N_A_M1010_g N_VPWR_c_838_n 0.00527225f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_261 N_A_c_163_n N_VPWR_c_839_n 0.00402941f $X=2.845 $Y=2.55 $X2=0 $Y2=0
cc_262 N_A_c_164_n N_VPWR_c_839_n 3.72682e-19 $X=3.265 $Y=2.475 $X2=0 $Y2=0
cc_263 N_A_c_167_n N_VPWR_c_839_n 0.00796123f $X=3.415 $Y=3.15 $X2=0 $Y2=0
cc_264 N_A_c_166_n N_VPWR_c_840_n 0.0188328f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_265 N_A_c_166_n N_VPWR_c_841_n 0.0676295f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_266 N_A_M1010_g N_VPWR_c_831_n 0.00975732f $X=1.015 $Y=2.87 $X2=0 $Y2=0
cc_267 N_A_c_163_n N_VPWR_c_831_n 0.00492937f $X=2.845 $Y=2.55 $X2=0 $Y2=0
cc_268 N_A_c_166_n N_VPWR_c_831_n 0.0238174f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_269 N_A_c_167_n N_VPWR_c_831_n 0.0103159f $X=3.415 $Y=3.15 $X2=0 $Y2=0
cc_270 N_A_c_169_n N_VPWR_c_831_n 0.0796388f $X=6.585 $Y=3.15 $X2=0 $Y2=0
cc_271 N_A_c_172_n N_VPWR_c_831_n 0.00888046f $X=4.79 $Y=3.15 $X2=0 $Y2=0
cc_272 N_A_c_163_n N_A_404_532#_c_928_n 0.00766076f $X=2.845 $Y=2.55 $X2=0 $Y2=0
cc_273 N_A_c_164_n N_A_404_532#_c_928_n 0.00829766f $X=3.265 $Y=2.475 $X2=0
+ $Y2=0
cc_274 N_A_c_165_n N_A_404_532#_c_928_n 0.00117858f $X=3.34 $Y=3.075 $X2=0 $Y2=0
cc_275 N_A_c_171_n N_A_404_532#_c_928_n 0.00367188f $X=2.845 $Y=2.475 $X2=0
+ $Y2=0
cc_276 N_A_c_165_n N_A_404_532#_c_930_n 0.0036237f $X=3.34 $Y=3.075 $X2=0 $Y2=0
cc_277 N_A_c_166_n N_A_781_457#_c_956_n 0.00444435f $X=4.715 $Y=3.15 $X2=0 $Y2=0
cc_278 N_A_M1013_g N_A_781_457#_c_956_n 3.54034e-19 $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_279 N_A_M1013_g N_A_781_457#_c_957_n 0.0151632f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_280 N_A_M1013_g N_A_781_457#_c_959_n 0.00561315f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_281 N_A_c_169_n N_A_781_457#_c_959_n 0.00321277f $X=6.585 $Y=3.15 $X2=0 $Y2=0
cc_282 N_A_M1003_g N_VGND_c_1004_n 0.0090565f $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_283 N_A_M1023_g N_VGND_c_1005_n 0.00453764f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_284 N_A_M1023_g N_VGND_c_1006_n 0.0041494f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_285 N_A_M1013_g N_VGND_c_1007_n 0.00381005f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_286 N_A_M1001_g N_VGND_c_1008_n 0.0173317f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_287 N_A_M1001_g N_VGND_c_1009_n 0.00429645f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_288 N_A_M1003_g N_VGND_c_1015_n 7.88961e-19 $X=1.045 $Y=0.805 $X2=0 $Y2=0
cc_289 N_A_M1023_g N_VGND_c_1015_n 9.39239e-19 $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_290 N_A_M1013_g N_VGND_c_1015_n 9.39239e-19 $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_291 N_A_M1001_g N_VGND_c_1015_n 0.00497858f $X=6.64 $Y=0.515 $X2=0 $Y2=0
cc_292 N_A_M1023_g N_A_382_119#_c_1096_n 0.00972361f $X=2.855 $Y=0.805 $X2=0
+ $Y2=0
cc_293 N_A_M1023_g N_A_382_119#_c_1097_n 6.19371e-19 $X=2.855 $Y=0.805 $X2=0
+ $Y2=0
cc_294 N_A_M1023_g N_A_382_119#_c_1098_n 0.00645993f $X=2.855 $Y=0.805 $X2=0
+ $Y2=0
cc_295 N_A_M1013_g N_A_781_119#_c_1125_n 3.76938e-19 $X=4.79 $Y=0.805 $X2=0
+ $Y2=0
cc_296 N_A_M1013_g N_A_781_119#_c_1123_n 0.014626f $X=4.79 $Y=0.805 $X2=0 $Y2=0
cc_297 N_A_M1013_g N_A_781_119#_c_1127_n 0.00543534f $X=4.79 $Y=0.805 $X2=0
+ $Y2=0
cc_298 N_B_M1020_g N_CIN_M1022_g 0.0135233f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_299 N_B_c_329_n N_CIN_M1022_g 0.0118624f $X=2.32 $Y=1.125 $X2=0 $Y2=0
cc_300 N_B_M1020_g N_CIN_M1005_g 0.0169469f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_301 N_B_M1025_g N_CIN_M1005_g 0.0216664f $X=1.405 $Y=2.87 $X2=0 $Y2=0
cc_302 N_B_M1021_g N_CIN_M1005_g 0.0200136f $X=2.375 $Y=2.87 $X2=0 $Y2=0
cc_303 N_B_c_340_n N_CIN_M1005_g 0.0190393f $X=3.13 $Y=2.155 $X2=0 $Y2=0
cc_304 N_B_c_341_n N_CIN_M1005_g 0.021335f $X=1.495 $Y=2.155 $X2=0 $Y2=0
cc_305 N_B_c_342_n N_CIN_M1005_g 0.021772f $X=2.395 $Y=2.235 $X2=0 $Y2=0
cc_306 N_B_M1017_g N_CIN_M1002_g 0.0366651f $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_307 N_B_M1018_g N_CIN_M1004_g 0.0187031f $X=4.26 $Y=2.495 $X2=0 $Y2=0
cc_308 N_B_c_343_n N_CIN_M1004_g 0.0164814f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_309 N_B_c_344_n N_CIN_M1004_g 0.0192649f $X=4.31 $Y=1.84 $X2=0 $Y2=0
cc_310 N_B_c_345_n N_CIN_M1004_g 0.00817597f $X=3.215 $Y=1.84 $X2=0 $Y2=0
cc_311 N_B_M1014_g N_CIN_M1012_g 0.0343727f $X=6.12 $Y=0.805 $X2=0 $Y2=0
cc_312 B N_CIN_M1012_g 5.41588e-19 $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_313 N_B_c_328_n N_CIN_M1019_g 0.0661688f $X=6.12 $Y=2.125 $X2=0 $Y2=0
cc_314 N_B_c_343_n N_CIN_M1019_g 0.016343f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_315 B N_CIN_M1019_g 6.96917e-19 $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_316 N_B_M1020_g N_CIN_c_496_n 7.60334e-19 $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_317 N_B_c_330_n N_CIN_c_496_n 0.00456235f $X=2.32 $Y=1.275 $X2=0 $Y2=0
cc_318 N_B_c_340_n N_CIN_c_496_n 0.00601162f $X=3.13 $Y=2.155 $X2=0 $Y2=0
cc_319 N_B_c_343_n N_CIN_c_496_n 0.00608749f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_320 N_B_c_345_n N_CIN_c_496_n 0.00838045f $X=3.215 $Y=1.84 $X2=0 $Y2=0
cc_321 N_B_c_332_n N_CIN_c_496_n 0.00682565f $X=2.395 $Y=2.07 $X2=0 $Y2=0
cc_322 N_B_M1020_g N_CIN_c_497_n 0.021044f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_323 N_B_c_330_n N_CIN_c_497_n 0.00860136f $X=2.32 $Y=1.275 $X2=0 $Y2=0
cc_324 N_B_c_332_n N_CIN_c_497_n 0.0449429f $X=2.395 $Y=2.07 $X2=0 $Y2=0
cc_325 N_B_M1014_g N_CIN_c_498_n 9.2777e-19 $X=6.12 $Y=0.805 $X2=0 $Y2=0
cc_326 B N_CIN_c_498_n 0.015117f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_327 N_B_M1014_g N_CIN_c_499_n 0.0198423f $X=6.12 $Y=0.805 $X2=0 $Y2=0
cc_328 N_B_c_343_n N_CIN_c_499_n 0.00455934f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_329 B N_CIN_c_499_n 5.59493e-19 $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_330 N_B_M1017_g N_CIN_c_500_n 0.0129954f $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_331 N_B_c_343_n N_CIN_c_500_n 0.150637f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_332 N_B_c_344_n N_CIN_c_500_n 0.00446495f $X=4.31 $Y=1.84 $X2=0 $Y2=0
cc_333 N_B_M1017_g N_CIN_c_501_n 8.85232e-19 $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_334 N_B_c_343_n N_CIN_c_501_n 0.028703f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_335 N_B_c_343_n N_CIN_c_502_n 0.00199112f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_336 N_B_M1020_g N_A_80_225#_c_612_n 0.00979198f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_337 N_B_M1017_g N_A_80_225#_c_612_n 0.0104164f $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_338 N_B_c_329_n N_A_80_225#_c_612_n 0.0100733f $X=2.32 $Y=1.125 $X2=0 $Y2=0
cc_339 N_B_c_343_n N_A_80_225#_M1024_g 0.0154085f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_340 N_B_M1020_g N_A_80_225#_c_618_n 0.00712331f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_341 N_B_c_340_n N_A_80_225#_c_625_n 0.0110795f $X=3.13 $Y=2.155 $X2=0 $Y2=0
cc_342 N_B_c_341_n N_A_80_225#_c_625_n 0.0022724f $X=1.495 $Y=2.155 $X2=0 $Y2=0
cc_343 N_B_M1025_g N_A_80_225#_c_627_n 0.00746098f $X=1.405 $Y=2.87 $X2=0 $Y2=0
cc_344 N_B_M1025_g N_A_80_225#_c_667_n 0.0189871f $X=1.405 $Y=2.87 $X2=0 $Y2=0
cc_345 N_B_c_340_n N_A_80_225#_c_667_n 0.016581f $X=3.13 $Y=2.155 $X2=0 $Y2=0
cc_346 N_B_c_341_n N_A_80_225#_c_667_n 0.0033386f $X=1.495 $Y=2.155 $X2=0 $Y2=0
cc_347 N_B_M1020_g N_A_80_225#_c_619_n 0.0041375f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_348 N_B_M1020_g N_A_80_225#_c_657_n 0.00861766f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_349 N_B_M1014_g N_A_1059_119#_c_741_n 0.0154129f $X=6.12 $Y=0.805 $X2=0 $Y2=0
cc_350 B N_A_1059_119#_c_741_n 0.0373057f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_351 N_B_c_328_n N_A_1059_119#_c_754_n 0.00114275f $X=6.12 $Y=2.125 $X2=0
+ $Y2=0
cc_352 N_B_M1009_g N_A_1059_119#_c_754_n 0.0115003f $X=6.12 $Y=2.495 $X2=0 $Y2=0
cc_353 N_B_c_343_n N_A_1059_119#_c_754_n 0.0522646f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_354 B N_A_1059_119#_c_742_n 0.0750525f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_355 N_B_M1014_g N_A_1059_119#_c_743_n 0.00107358f $X=6.12 $Y=0.805 $X2=0
+ $Y2=0
cc_356 N_B_c_343_n N_A_1059_119#_c_759_n 0.0129093f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_357 N_B_M1021_g N_VPWR_c_833_n 0.00679722f $X=2.375 $Y=2.87 $X2=0 $Y2=0
cc_358 N_B_c_343_n N_VPWR_c_834_n 0.0111515f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_359 N_B_M1018_g N_VPWR_c_835_n 0.00207537f $X=4.26 $Y=2.495 $X2=0 $Y2=0
cc_360 N_B_M1025_g N_VPWR_c_838_n 0.00355856f $X=1.405 $Y=2.87 $X2=0 $Y2=0
cc_361 N_B_M1021_g N_VPWR_c_838_n 0.00402941f $X=2.375 $Y=2.87 $X2=0 $Y2=0
cc_362 N_B_M1025_g N_VPWR_c_831_n 0.00545466f $X=1.405 $Y=2.87 $X2=0 $Y2=0
cc_363 N_B_M1021_g N_VPWR_c_831_n 0.00480023f $X=2.375 $Y=2.87 $X2=0 $Y2=0
cc_364 N_B_M1018_g N_VPWR_c_831_n 9.49986e-19 $X=4.26 $Y=2.495 $X2=0 $Y2=0
cc_365 N_B_M1009_g N_VPWR_c_831_n 9.49986e-19 $X=6.12 $Y=2.495 $X2=0 $Y2=0
cc_366 N_B_M1025_g N_A_404_532#_c_936_n 4.33604e-19 $X=1.405 $Y=2.87 $X2=0 $Y2=0
cc_367 N_B_M1021_g N_A_404_532#_c_928_n 0.0120148f $X=2.375 $Y=2.87 $X2=0 $Y2=0
cc_368 N_B_c_340_n N_A_404_532#_c_928_n 0.0652668f $X=3.13 $Y=2.155 $X2=0 $Y2=0
cc_369 N_B_c_342_n N_A_404_532#_c_928_n 0.00343224f $X=2.395 $Y=2.235 $X2=0
+ $Y2=0
cc_370 N_B_c_345_n N_A_404_532#_c_928_n 0.0081283f $X=3.215 $Y=1.84 $X2=0 $Y2=0
cc_371 N_B_M1025_g N_A_404_532#_c_929_n 7.81771e-19 $X=1.405 $Y=2.87 $X2=0 $Y2=0
cc_372 N_B_c_340_n N_A_404_532#_c_929_n 0.0239459f $X=3.13 $Y=2.155 $X2=0 $Y2=0
cc_373 N_B_c_342_n N_A_404_532#_c_929_n 0.00121025f $X=2.395 $Y=2.235 $X2=0
+ $Y2=0
cc_374 N_B_M1018_g N_A_781_457#_c_956_n 0.00560651f $X=4.26 $Y=2.495 $X2=0 $Y2=0
cc_375 N_B_c_345_n N_A_781_457#_c_956_n 0.00113648f $X=3.215 $Y=1.84 $X2=0 $Y2=0
cc_376 N_B_M1018_g N_A_781_457#_c_957_n 0.0128172f $X=4.26 $Y=2.495 $X2=0 $Y2=0
cc_377 N_B_c_343_n N_A_781_457#_c_957_n 0.0713576f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_378 N_B_c_344_n N_A_781_457#_c_957_n 0.00345061f $X=4.31 $Y=1.84 $X2=0 $Y2=0
cc_379 N_B_M1018_g N_A_781_457#_c_958_n 0.00176361f $X=4.26 $Y=2.495 $X2=0 $Y2=0
cc_380 N_B_c_343_n N_A_781_457#_c_958_n 0.0227007f $X=6.01 $Y=1.84 $X2=0 $Y2=0
cc_381 N_B_c_344_n N_A_781_457#_c_958_n 0.00101959f $X=4.31 $Y=1.84 $X2=0 $Y2=0
cc_382 N_B_c_345_n N_A_781_457#_c_958_n 0.00578528f $X=3.215 $Y=1.84 $X2=0 $Y2=0
cc_383 N_B_M1018_g N_A_781_457#_c_959_n 3.53882e-19 $X=4.26 $Y=2.495 $X2=0 $Y2=0
cc_384 N_B_M1020_g N_VGND_c_1004_n 0.00117548f $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_385 N_B_c_329_n N_VGND_c_1005_n 0.00453764f $X=2.32 $Y=1.125 $X2=0 $Y2=0
cc_386 N_B_M1017_g N_VGND_c_1006_n 4.3095e-19 $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_387 N_B_M1017_g N_VGND_c_1007_n 0.00201884f $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_388 N_B_M1014_g N_VGND_c_1008_n 0.00100768f $X=6.12 $Y=0.805 $X2=0 $Y2=0
cc_389 N_B_M1014_g N_VGND_c_1009_n 0.00431487f $X=6.12 $Y=0.805 $X2=0 $Y2=0
cc_390 N_B_M1020_g N_VGND_c_1015_n 9.39239e-19 $X=1.405 $Y=0.805 $X2=0 $Y2=0
cc_391 N_B_M1017_g N_VGND_c_1015_n 9.39239e-19 $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_392 N_B_M1014_g N_VGND_c_1015_n 0.00477801f $X=6.12 $Y=0.805 $X2=0 $Y2=0
cc_393 N_B_c_329_n N_VGND_c_1015_n 9.39239e-19 $X=2.32 $Y=1.125 $X2=0 $Y2=0
cc_394 N_B_c_329_n N_A_382_119#_c_1096_n 0.00969482f $X=2.32 $Y=1.125 $X2=0
+ $Y2=0
cc_395 N_B_c_330_n N_A_382_119#_c_1096_n 8.94506e-19 $X=2.32 $Y=1.275 $X2=0
+ $Y2=0
cc_396 N_B_c_329_n N_A_382_119#_c_1097_n 0.00594029f $X=2.32 $Y=1.125 $X2=0
+ $Y2=0
cc_397 N_B_c_329_n N_A_382_119#_c_1098_n 6.19475e-19 $X=2.32 $Y=1.125 $X2=0
+ $Y2=0
cc_398 N_B_M1017_g N_A_781_119#_c_1125_n 0.00548392f $X=4.26 $Y=0.805 $X2=0
+ $Y2=0
cc_399 N_B_M1017_g N_A_781_119#_c_1123_n 0.0128075f $X=4.26 $Y=0.805 $X2=0 $Y2=0
cc_400 N_B_M1017_g N_A_781_119#_c_1124_n 0.00162261f $X=4.26 $Y=0.805 $X2=0
+ $Y2=0
cc_401 N_B_M1017_g N_A_781_119#_c_1127_n 3.76105e-19 $X=4.26 $Y=0.805 $X2=0
+ $Y2=0
cc_402 N_CIN_M1022_g N_A_80_225#_c_612_n 0.0104164f $X=1.835 $Y=0.805 $X2=0
+ $Y2=0
cc_403 N_CIN_M1002_g N_A_80_225#_c_612_n 0.0103107f $X=3.83 $Y=0.805 $X2=0 $Y2=0
cc_404 N_CIN_M1012_g N_A_80_225#_M1011_g 0.0211972f $X=5.65 $Y=0.805 $X2=0 $Y2=0
cc_405 N_CIN_M1019_g N_A_80_225#_M1024_g 0.0306584f $X=5.73 $Y=2.495 $X2=0 $Y2=0
cc_406 N_CIN_c_498_n N_A_80_225#_M1024_g 4.61159e-19 $X=5.67 $Y=1.46 $X2=0 $Y2=0
cc_407 N_CIN_c_499_n N_A_80_225#_M1024_g 0.0212031f $X=5.67 $Y=1.46 $X2=0 $Y2=0
cc_408 N_CIN_c_500_n N_A_80_225#_M1024_g 0.0164872f $X=5.505 $Y=1.44 $X2=0 $Y2=0
cc_409 N_CIN_c_500_n N_A_80_225#_c_616_n 7.21492e-19 $X=5.505 $Y=1.44 $X2=0
+ $Y2=0
cc_410 N_CIN_M1022_g N_A_80_225#_c_618_n 6.312e-19 $X=1.835 $Y=0.805 $X2=0 $Y2=0
cc_411 N_CIN_c_496_n N_A_80_225#_c_618_n 0.00570588f $X=3.435 $Y=1.315 $X2=0
+ $Y2=0
cc_412 N_CIN_c_497_n N_A_80_225#_c_618_n 0.00245112f $X=1.855 $Y=1.315 $X2=0
+ $Y2=0
cc_413 N_CIN_M1022_g N_A_80_225#_c_619_n 0.00170372f $X=1.835 $Y=0.805 $X2=0
+ $Y2=0
cc_414 N_CIN_c_496_n N_A_80_225#_c_657_n 0.00170864f $X=3.435 $Y=1.315 $X2=0
+ $Y2=0
cc_415 N_CIN_c_497_n N_A_80_225#_c_657_n 0.00114847f $X=1.855 $Y=1.315 $X2=0
+ $Y2=0
cc_416 N_CIN_M1012_g N_A_1059_119#_c_741_n 0.0100453f $X=5.65 $Y=0.805 $X2=0
+ $Y2=0
cc_417 N_CIN_c_498_n N_A_1059_119#_c_741_n 0.01181f $X=5.67 $Y=1.46 $X2=0 $Y2=0
cc_418 N_CIN_c_499_n N_A_1059_119#_c_741_n 0.00258162f $X=5.67 $Y=1.46 $X2=0
+ $Y2=0
cc_419 N_CIN_M1019_g N_A_1059_119#_c_754_n 0.0100793f $X=5.73 $Y=2.495 $X2=0
+ $Y2=0
cc_420 N_CIN_M1012_g N_A_1059_119#_c_743_n 0.00589191f $X=5.65 $Y=0.805 $X2=0
+ $Y2=0
cc_421 N_CIN_c_498_n N_A_1059_119#_c_743_n 0.00513822f $X=5.67 $Y=1.46 $X2=0
+ $Y2=0
cc_422 N_CIN_c_499_n N_A_1059_119#_c_743_n 0.00150197f $X=5.67 $Y=1.46 $X2=0
+ $Y2=0
cc_423 N_CIN_c_500_n N_A_1059_119#_c_743_n 0.00973267f $X=5.505 $Y=1.44 $X2=0
+ $Y2=0
cc_424 N_CIN_M1005_g N_VPWR_c_833_n 0.00109992f $X=1.945 $Y=2.87 $X2=0 $Y2=0
cc_425 N_CIN_M1004_g N_VPWR_c_834_n 0.00212242f $X=3.83 $Y=2.495 $X2=0 $Y2=0
cc_426 N_CIN_M1005_g N_VPWR_c_838_n 0.00535803f $X=1.945 $Y=2.87 $X2=0 $Y2=0
cc_427 N_CIN_M1005_g N_VPWR_c_831_n 0.01021f $X=1.945 $Y=2.87 $X2=0 $Y2=0
cc_428 N_CIN_M1004_g N_VPWR_c_831_n 9.49986e-19 $X=3.83 $Y=2.495 $X2=0 $Y2=0
cc_429 N_CIN_M1019_g N_VPWR_c_831_n 9.49986e-19 $X=5.73 $Y=2.495 $X2=0 $Y2=0
cc_430 N_CIN_M1005_g N_A_404_532#_c_936_n 0.00461209f $X=1.945 $Y=2.87 $X2=0
+ $Y2=0
cc_431 N_CIN_M1005_g N_A_404_532#_c_929_n 0.00599561f $X=1.945 $Y=2.87 $X2=0
+ $Y2=0
cc_432 N_CIN_M1004_g N_A_781_457#_c_956_n 3.66692e-19 $X=3.83 $Y=2.495 $X2=0
+ $Y2=0
cc_433 N_CIN_M1019_g N_A_781_457#_c_957_n 7.59826e-19 $X=5.73 $Y=2.495 $X2=0
+ $Y2=0
cc_434 N_CIN_M1004_g N_A_781_457#_c_958_n 0.00293045f $X=3.83 $Y=2.495 $X2=0
+ $Y2=0
cc_435 N_CIN_M1002_g N_VGND_c_1006_n 0.00971164f $X=3.83 $Y=0.805 $X2=0 $Y2=0
cc_436 N_CIN_c_501_n N_VGND_c_1006_n 0.0265395f $X=3.6 $Y=1.375 $X2=0 $Y2=0
cc_437 N_CIN_c_502_n N_VGND_c_1006_n 0.00180983f $X=3.83 $Y=1.375 $X2=0 $Y2=0
cc_438 N_CIN_M1012_g N_VGND_c_1009_n 0.00415648f $X=5.65 $Y=0.805 $X2=0 $Y2=0
cc_439 N_CIN_M1022_g N_VGND_c_1015_n 9.39239e-19 $X=1.835 $Y=0.805 $X2=0 $Y2=0
cc_440 N_CIN_M1002_g N_VGND_c_1015_n 7.88961e-19 $X=3.83 $Y=0.805 $X2=0 $Y2=0
cc_441 N_CIN_M1012_g N_VGND_c_1015_n 0.00477801f $X=5.65 $Y=0.805 $X2=0 $Y2=0
cc_442 N_CIN_c_496_n N_A_382_119#_c_1096_n 0.0483073f $X=3.435 $Y=1.315 $X2=0
+ $Y2=0
cc_443 N_CIN_M1022_g N_A_382_119#_c_1097_n 6.45781e-19 $X=1.835 $Y=0.805 $X2=0
+ $Y2=0
cc_444 N_CIN_c_496_n N_A_382_119#_c_1097_n 0.0261281f $X=3.435 $Y=1.315 $X2=0
+ $Y2=0
cc_445 N_CIN_c_497_n N_A_382_119#_c_1097_n 0.00307463f $X=1.855 $Y=1.315 $X2=0
+ $Y2=0
cc_446 N_CIN_M1002_g N_A_382_119#_c_1098_n 0.00221061f $X=3.83 $Y=0.805 $X2=0
+ $Y2=0
cc_447 N_CIN_c_496_n N_A_382_119#_c_1098_n 0.0257096f $X=3.435 $Y=1.315 $X2=0
+ $Y2=0
cc_448 N_CIN_M1002_g N_A_781_119#_c_1125_n 3.15901e-19 $X=3.83 $Y=0.805 $X2=0
+ $Y2=0
cc_449 N_CIN_M1012_g N_A_781_119#_c_1123_n 3.20072e-19 $X=5.65 $Y=0.805 $X2=0
+ $Y2=0
cc_450 N_CIN_c_500_n N_A_781_119#_c_1123_n 0.0727345f $X=5.505 $Y=1.44 $X2=0
+ $Y2=0
cc_451 N_CIN_M1002_g N_A_781_119#_c_1124_n 0.00384623f $X=3.83 $Y=0.805 $X2=0
+ $Y2=0
cc_452 N_CIN_c_500_n N_A_781_119#_c_1124_n 0.0194394f $X=5.505 $Y=1.44 $X2=0
+ $Y2=0
cc_453 N_CIN_c_501_n N_A_781_119#_c_1124_n 0.00551883f $X=3.6 $Y=1.375 $X2=0
+ $Y2=0
cc_454 N_A_80_225#_c_621_n N_COUT_c_814_n 0.00397231f $X=0.59 $Y=1.29 $X2=0
+ $Y2=0
cc_455 N_A_80_225#_M1007_g N_COUT_c_816_n 0.00876323f $X=0.475 $Y=2.76 $X2=0
+ $Y2=0
cc_456 N_A_80_225#_c_627_n N_COUT_c_816_n 0.00382731f $X=1.145 $Y=2.705 $X2=0
+ $Y2=0
cc_457 N_A_80_225#_M1026_g COUT 0.00527823f $X=0.615 $Y=0.805 $X2=0 $Y2=0
cc_458 N_A_80_225#_c_617_n COUT 0.0472521f $X=0.615 $Y=2.195 $X2=0 $Y2=0
cc_459 N_A_80_225#_c_626_n COUT 0.012116f $X=0.7 $Y=2.28 $X2=0 $Y2=0
cc_460 N_A_80_225#_c_620_n COUT 0.0245945f $X=0.597 $Y=1.21 $X2=0 $Y2=0
cc_461 N_A_80_225#_c_621_n COUT 0.0328169f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_462 N_A_80_225#_M1007_g N_VPWR_c_832_n 0.00335592f $X=0.475 $Y=2.76 $X2=0
+ $Y2=0
cc_463 N_A_80_225#_c_625_n N_VPWR_c_832_n 0.0103069f $X=1.06 $Y=2.28 $X2=0 $Y2=0
cc_464 N_A_80_225#_c_626_n N_VPWR_c_832_n 0.00606502f $X=0.7 $Y=2.28 $X2=0 $Y2=0
cc_465 N_A_80_225#_M1007_g N_VPWR_c_837_n 0.00534537f $X=0.475 $Y=2.76 $X2=0
+ $Y2=0
cc_466 N_A_80_225#_c_653_n N_VPWR_c_838_n 0.0078668f $X=1.23 $Y=2.87 $X2=0 $Y2=0
cc_467 N_A_80_225#_c_667_n N_VPWR_c_838_n 0.0280814f $X=1.685 $Y=2.87 $X2=0
+ $Y2=0
cc_468 N_A_80_225#_M1007_g N_VPWR_c_831_n 0.0109328f $X=0.475 $Y=2.76 $X2=0
+ $Y2=0
cc_469 N_A_80_225#_M1024_g N_VPWR_c_831_n 9.49986e-19 $X=5.22 $Y=2.495 $X2=0
+ $Y2=0
cc_470 N_A_80_225#_c_653_n N_VPWR_c_831_n 0.00633145f $X=1.23 $Y=2.87 $X2=0
+ $Y2=0
cc_471 N_A_80_225#_c_667_n N_VPWR_c_831_n 0.0214901f $X=1.685 $Y=2.87 $X2=0
+ $Y2=0
cc_472 N_A_80_225#_c_627_n A_218_532# 4.90897e-19 $X=1.145 $Y=2.705 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_80_225#_c_653_n A_218_532# 8.73591e-19 $X=1.23 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_474 N_A_80_225#_c_667_n A_218_532# 0.00217459f $X=1.685 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_475 N_A_80_225#_M1024_g N_A_781_457#_c_957_n 0.00575952f $X=5.22 $Y=2.495
+ $X2=0 $Y2=0
cc_476 N_A_80_225#_M1024_g N_A_781_457#_c_959_n 6.12464e-19 $X=5.22 $Y=2.495
+ $X2=0 $Y2=0
cc_477 N_A_80_225#_M1026_g N_VGND_c_1004_n 0.0258004f $X=0.615 $Y=0.805 $X2=0
+ $Y2=0
cc_478 N_A_80_225#_c_612_n N_VGND_c_1004_n 0.0183562f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_479 N_A_80_225#_c_613_n N_VGND_c_1004_n 0.00388727f $X=0.69 $Y=0.18 $X2=0
+ $Y2=0
cc_480 N_A_80_225#_c_618_n N_VGND_c_1004_n 0.0192379f $X=1.255 $Y=1.21 $X2=0
+ $Y2=0
cc_481 N_A_80_225#_c_620_n N_VGND_c_1004_n 0.00237022f $X=0.597 $Y=1.21 $X2=0
+ $Y2=0
cc_482 N_A_80_225#_c_621_n N_VGND_c_1004_n 0.0011583f $X=0.59 $Y=1.29 $X2=0
+ $Y2=0
cc_483 N_A_80_225#_c_657_n N_VGND_c_1004_n 0.0182155f $X=1.62 $Y=0.805 $X2=0
+ $Y2=0
cc_484 N_A_80_225#_c_612_n N_VGND_c_1005_n 0.0255378f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_485 N_A_80_225#_c_612_n N_VGND_c_1006_n 0.0247996f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_486 N_A_80_225#_c_612_n N_VGND_c_1007_n 0.0248734f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_487 N_A_80_225#_M1011_g N_VGND_c_1007_n 0.00602502f $X=5.22 $Y=0.805 $X2=0
+ $Y2=0
cc_488 N_A_80_225#_c_612_n N_VGND_c_1009_n 0.019224f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_489 N_A_80_225#_c_612_n N_VGND_c_1011_n 0.0413845f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_490 N_A_80_225#_c_657_n N_VGND_c_1011_n 0.00734684f $X=1.62 $Y=0.805 $X2=0
+ $Y2=0
cc_491 N_A_80_225#_c_612_n N_VGND_c_1012_n 0.0214644f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_492 N_A_80_225#_c_612_n N_VGND_c_1013_n 0.0179878f $X=5.145 $Y=0.18 $X2=0
+ $Y2=0
cc_493 N_A_80_225#_c_612_n N_VGND_c_1015_n 0.11565f $X=5.145 $Y=0.18 $X2=0 $Y2=0
cc_494 N_A_80_225#_c_613_n N_VGND_c_1015_n 0.00947588f $X=0.69 $Y=0.18 $X2=0
+ $Y2=0
cc_495 N_A_80_225#_c_657_n N_VGND_c_1015_n 0.0122191f $X=1.62 $Y=0.805 $X2=0
+ $Y2=0
cc_496 N_A_80_225#_c_613_n N_VGND_c_1016_n 0.00486043f $X=0.69 $Y=0.18 $X2=0
+ $Y2=0
cc_497 N_A_80_225#_c_619_n A_224_119# 5.89303e-19 $X=1.387 $Y=1.125 $X2=-0.19
+ $Y2=-0.245
cc_498 N_A_80_225#_c_657_n A_224_119# 0.00366513f $X=1.62 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_499 N_A_80_225#_c_612_n N_A_382_119#_c_1096_n 0.00168455f $X=5.145 $Y=0.18
+ $X2=0 $Y2=0
cc_500 N_A_80_225#_c_612_n N_A_382_119#_c_1097_n 0.00532861f $X=5.145 $Y=0.18
+ $X2=0 $Y2=0
cc_501 N_A_80_225#_c_619_n N_A_382_119#_c_1097_n 0.00200432f $X=1.387 $Y=1.125
+ $X2=0 $Y2=0
cc_502 N_A_80_225#_c_612_n N_A_382_119#_c_1098_n 0.00540587f $X=5.145 $Y=0.18
+ $X2=0 $Y2=0
cc_503 N_A_80_225#_c_612_n N_A_781_119#_c_1125_n 0.00396815f $X=5.145 $Y=0.18
+ $X2=0 $Y2=0
cc_504 N_A_80_225#_M1011_g N_A_781_119#_c_1123_n 0.00336213f $X=5.22 $Y=0.805
+ $X2=0 $Y2=0
cc_505 N_A_80_225#_c_616_n N_A_781_119#_c_1123_n 0.00288973f $X=5.205 $Y=1.275
+ $X2=0 $Y2=0
cc_506 N_A_80_225#_c_612_n N_A_781_119#_c_1127_n 0.00332259f $X=5.145 $Y=0.18
+ $X2=0 $Y2=0
cc_507 N_A_80_225#_M1011_g N_A_781_119#_c_1127_n 2.70691e-19 $X=5.22 $Y=0.805
+ $X2=0 $Y2=0
cc_508 N_A_1059_119#_c_754_n N_VPWR_M1015_d 0.00433709f $X=6.745 $Y=2.38 $X2=0
+ $Y2=0
cc_509 N_A_1059_119#_M1000_g N_VPWR_c_836_n 0.00917425f $X=7.205 $Y=2.605 $X2=0
+ $Y2=0
cc_510 N_A_1059_119#_c_754_n N_VPWR_c_836_n 0.0130971f $X=6.745 $Y=2.38 $X2=0
+ $Y2=0
cc_511 N_A_1059_119#_c_759_n N_VPWR_c_841_n 0.00499893f $X=5.48 $Y=2.38 $X2=0
+ $Y2=0
cc_512 N_A_1059_119#_M1000_g N_VPWR_c_842_n 0.00532616f $X=7.205 $Y=2.605 $X2=0
+ $Y2=0
cc_513 N_A_1059_119#_M1000_g N_VPWR_c_831_n 0.00520409f $X=7.205 $Y=2.605 $X2=0
+ $Y2=0
cc_514 N_A_1059_119#_c_754_n N_VPWR_c_831_n 0.00285456f $X=6.745 $Y=2.38 $X2=0
+ $Y2=0
cc_515 N_A_1059_119#_c_759_n N_VPWR_c_831_n 0.00818309f $X=5.48 $Y=2.38 $X2=0
+ $Y2=0
cc_516 N_A_1059_119#_c_754_n A_1161_457# 0.00407027f $X=6.745 $Y=2.38 $X2=-0.19
+ $Y2=-0.245
cc_517 N_A_1059_119#_c_754_n A_1239_457# 0.00828386f $X=6.745 $Y=2.38 $X2=-0.19
+ $Y2=-0.245
cc_518 N_A_1059_119#_c_747_n N_SUM_c_987_n 0.00467152f $X=7.09 $Y=1.03 $X2=0
+ $Y2=0
cc_519 N_A_1059_119#_M1000_g N_SUM_c_988_n 0.0234449f $X=7.205 $Y=2.605 $X2=0
+ $Y2=0
cc_520 N_A_1059_119#_c_742_n N_SUM_c_988_n 0.0425707f $X=6.85 $Y=2.295 $X2=0
+ $Y2=0
cc_521 N_A_1059_119#_c_742_n SUM 0.00925956f $X=6.85 $Y=2.295 $X2=0 $Y2=0
cc_522 N_A_1059_119#_c_746_n SUM 0.0276957f $X=7.09 $Y=1.03 $X2=0 $Y2=0
cc_523 N_A_1059_119#_c_747_n SUM 0.0149279f $X=7.09 $Y=1.03 $X2=0 $Y2=0
cc_524 N_A_1059_119#_c_748_n SUM 0.00487247f $X=7.102 $Y=0.835 $X2=0 $Y2=0
cc_525 N_A_1059_119#_c_745_n N_VGND_c_1008_n 0.0195971f $X=6.745 $Y=1.022 $X2=0
+ $Y2=0
cc_526 N_A_1059_119#_c_747_n N_VGND_c_1008_n 0.00127937f $X=7.09 $Y=1.03 $X2=0
+ $Y2=0
cc_527 N_A_1059_119#_c_748_n N_VGND_c_1008_n 0.00337322f $X=7.102 $Y=0.835 $X2=0
+ $Y2=0
cc_528 N_A_1059_119#_c_743_n N_VGND_c_1009_n 0.00449519f $X=5.435 $Y=0.795 $X2=0
+ $Y2=0
cc_529 N_A_1059_119#_c_748_n N_VGND_c_1014_n 0.0051746f $X=7.102 $Y=0.835 $X2=0
+ $Y2=0
cc_530 N_A_1059_119#_c_741_n N_VGND_c_1015_n 0.0312164f $X=6.428 $Y=0.927 $X2=0
+ $Y2=0
cc_531 N_A_1059_119#_c_743_n N_VGND_c_1015_n 0.00851503f $X=5.435 $Y=0.795 $X2=0
+ $Y2=0
cc_532 N_A_1059_119#_c_745_n N_VGND_c_1015_n 0.00588864f $X=6.745 $Y=1.022 $X2=0
+ $Y2=0
cc_533 N_A_1059_119#_c_746_n N_VGND_c_1015_n 0.00508431f $X=7.09 $Y=1.03 $X2=0
+ $Y2=0
cc_534 N_A_1059_119#_c_747_n N_VGND_c_1015_n 5.10052e-19 $X=7.09 $Y=1.03 $X2=0
+ $Y2=0
cc_535 N_A_1059_119#_c_748_n N_VGND_c_1015_n 0.00611102f $X=7.102 $Y=0.835 $X2=0
+ $Y2=0
cc_536 N_A_1059_119#_c_743_n N_A_781_119#_c_1127_n 3.25523e-19 $X=5.435 $Y=0.795
+ $X2=0 $Y2=0
cc_537 N_A_1059_119#_c_741_n A_1145_119# 0.00416643f $X=6.428 $Y=0.927 $X2=-0.19
+ $Y2=-0.245
cc_538 N_A_1059_119#_c_741_n A_1239_119# 0.00363852f $X=6.428 $Y=0.927 $X2=-0.19
+ $Y2=-0.245
cc_539 N_A_1059_119#_c_744_n A_1239_119# 5.46085e-19 $X=6.52 $Y=0.927 $X2=-0.19
+ $Y2=-0.245
cc_540 N_COUT_c_816_n N_VPWR_c_837_n 0.0217292f $X=0.26 $Y=2.585 $X2=0 $Y2=0
cc_541 N_COUT_c_816_n N_VPWR_c_831_n 0.0130045f $X=0.26 $Y=2.585 $X2=0 $Y2=0
cc_542 N_COUT_c_814_n N_VGND_c_1015_n 0.0121257f $X=0.4 $Y=0.79 $X2=0 $Y2=0
cc_543 N_COUT_c_814_n N_VGND_c_1016_n 0.00771626f $X=0.4 $Y=0.79 $X2=0 $Y2=0
cc_544 N_VPWR_c_838_n N_A_404_532#_c_936_n 0.0129103f $X=2.445 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_831_n N_A_404_532#_c_936_n 0.0104015f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_833_n N_A_404_532#_c_928_n 0.0205348f $X=2.61 $Y=2.93 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_834_n N_A_404_532#_c_928_n 0.0111935f $X=3.615 $Y=2.49 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_838_n N_A_404_532#_c_928_n 0.00259279f $X=2.445 $Y=3.33 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_839_n N_A_404_532#_c_928_n 0.00259279f $X=3.47 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_831_n N_A_404_532#_c_928_n 0.0094343f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_834_n N_A_404_532#_c_930_n 0.0235063f $X=3.615 $Y=2.49 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_839_n N_A_404_532#_c_930_n 0.0145241f $X=3.47 $Y=3.33 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_831_n N_A_404_532#_c_930_n 0.0105246f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_840_n N_A_781_457#_c_956_n 0.00395476f $X=4.36 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_831_n N_A_781_457#_c_956_n 0.00694892f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_835_n N_A_781_457#_c_957_n 0.0243395f $X=4.525 $Y=2.54 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_841_n N_A_781_457#_c_959_n 0.00404585f $X=6.805 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_831_n N_A_781_457#_c_959_n 0.00718567f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_836_n SUM 0.0124071f $X=6.97 $Y=2.745 $X2=0 $Y2=0
cc_560 N_VPWR_c_842_n SUM 0.011264f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_561 N_VPWR_c_831_n SUM 0.0104094f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_562 N_SUM_c_987_n N_VGND_c_1014_n 0.0174397f $X=7.47 $Y=0.515 $X2=0 $Y2=0
cc_563 N_SUM_c_987_n N_VGND_c_1015_n 0.0158623f $X=7.47 $Y=0.515 $X2=0 $Y2=0
cc_564 N_VGND_M1027_d N_A_382_119#_c_1096_n 0.00307853f $X=2.38 $Y=0.595 $X2=0
+ $Y2=0
cc_565 N_VGND_c_1005_n N_A_382_119#_c_1096_n 0.0232685f $X=2.58 $Y=0.615 $X2=0
+ $Y2=0
cc_566 N_VGND_c_1011_n N_A_382_119#_c_1097_n 0.00507094f $X=2.415 $Y=0 $X2=0
+ $Y2=0
cc_567 N_VGND_c_1015_n N_A_382_119#_c_1097_n 0.00838363f $X=7.44 $Y=0 $X2=0
+ $Y2=0
cc_568 N_VGND_c_1006_n N_A_382_119#_c_1098_n 0.0225534f $X=3.615 $Y=0.795 $X2=0
+ $Y2=0
cc_569 N_VGND_c_1012_n N_A_382_119#_c_1098_n 0.00536621f $X=3.45 $Y=0 $X2=0
+ $Y2=0
cc_570 N_VGND_c_1015_n N_A_382_119#_c_1098_n 0.00812716f $X=7.44 $Y=0 $X2=0
+ $Y2=0
cc_571 N_VGND_c_1013_n N_A_781_119#_c_1125_n 0.00383003f $X=4.36 $Y=0 $X2=0
+ $Y2=0
cc_572 N_VGND_c_1015_n N_A_781_119#_c_1125_n 0.00596289f $X=7.44 $Y=0 $X2=0
+ $Y2=0
cc_573 N_VGND_c_1007_n N_A_781_119#_c_1123_n 0.0243395f $X=4.525 $Y=0.74 $X2=0
+ $Y2=0
cc_574 N_VGND_c_1009_n N_A_781_119#_c_1127_n 0.00432746f $X=6.69 $Y=0 $X2=0
+ $Y2=0
cc_575 N_VGND_c_1015_n N_A_781_119#_c_1127_n 0.00728309f $X=7.44 $Y=0 $X2=0
+ $Y2=0
