* File: sky130_fd_sc_lp__sdfxtp_lp.spice
* Created: Fri Aug 28 11:31:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfxtp_lp.pex.spice"
.subckt sky130_fd_sc_lp__sdfxtp_lp  VNB VPB D SCE SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* SCE	SCE
* D	D
* VPB	VPB
* VNB	VNB
MM1032 A_159_125# N_SCE_M1032_g N_A_27_409#_M1032_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_SCE_M1015_g A_159_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1025 A_351_125# N_A_27_409#_M1025_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=39.996 M=1 R=2.8 SA=75001.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_351_417#_M1003_d N_D_M1003_g A_351_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1034 A_531_125# N_SCE_M1034_g N_A_351_417#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0756 PD=0.73 PS=0.78 NRD=28.56 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_SCD_M1019_g A_531_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0651 PD=1.4 PS=0.73 NRD=0 NRS=28.56 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 A_820_66# N_CLK_M1018_g N_A_733_66#_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_CLK_M1020_g A_820_66# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1004 A_978_66# N_A_733_66#_M1004_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_A_998_347#_M1027_d N_A_733_66#_M1027_g A_978_66# VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_1263_155#_M1023_d N_A_998_347#_M1023_g N_A_1160_155#_M1023_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.1155 AS=0.1533 PD=0.97 PS=1.57 NRD=77.136 NRS=22.848
+ M=1 R=2.8 SA=75000.3 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1009 N_A_351_417#_M1009_d N_A_733_66#_M1009_g N_A_1263_155#_M1023_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1176 AS=0.1155 PD=1.4 PS=0.97 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_1576_99#_M1037_g N_A_1160_155#_M1037_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1211 AS=0.1197 PD=1.07 PS=1.41 NRD=66.66 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1028 A_1722_125# N_A_1263_155#_M1028_g N_VGND_M1037_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1211 PD=0.63 PS=1.07 NRD=14.28 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_A_1576_99#_M1016_d N_A_1263_155#_M1016_g A_1722_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_1957_347#_M1008_d N_A_733_66#_M1008_g N_A_1910_155#_M1008_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_1576_99#_M1010_d N_A_998_347#_M1010_g N_A_1957_347#_M1008_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.2521 AS=0.0588 PD=2.71 PS=0.7 NRD=155.772 NRS=0 M=1
+ R=2.8 SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_2148_185#_M1001_g N_A_1910_155#_M1001_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1024 A_2359_69# N_A_1957_347#_M1024_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_2148_185#_M1013_d N_A_1957_347#_M1013_g A_2359_69# VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_2628_69# N_A_2148_185#_M1002_g N_Q_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_2148_185#_M1035_g A_2628_69# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_SCE_M1005_g N_A_27_409#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.28 AS=0.285 PD=2.56 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1011 N_A_351_417#_M1011_d N_A_27_409#_M1011_g N_A_244_417#_M1011_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1000 A_457_417# N_D_M1000_g N_A_351_417#_M1011_d VPB PHIGHVT L=0.25 W=1
+ AD=0.11 AS=0.14 PD=1.22 PS=1.28 NRD=10.8153 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1030 N_VPWR_M1030_d N_SCE_M1030_g A_457_417# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.11 PD=1.28 PS=1.22 NRD=0 NRS=10.8153 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1014 N_A_244_417#_M1014_d N_SCD_M1014_g N_VPWR_M1030_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1029 N_VPWR_M1029_d N_CLK_M1029_g N_A_733_66#_M1029_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1012 N_A_998_347#_M1012_d N_A_733_66#_M1012_g N_VPWR_M1029_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1021 N_A_1263_155#_M1021_d N_A_998_347#_M1021_g N_A_351_417#_M1021_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4
+ SA=125000 SB=125005 A=0.25 P=2.5 MULT=1
MM1007 A_1528_347# N_A_733_66#_M1007_g N_A_1263_155#_M1021_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125001
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1022 N_VPWR_M1022_d N_A_1576_99#_M1022_g A_1528_347# VPB PHIGHVT L=0.25 W=1
+ AD=0.3525 AS=0.12 PD=1.705 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1036 N_A_1576_99#_M1036_d N_A_1263_155#_M1036_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.225 AS=0.3525 PD=1.45 PS=1.705 NRD=8.8453 NRS=83.7053 M=1 R=4
+ SA=125002 SB=125003 A=0.25 P=2.5 MULT=1
MM1017 N_A_1957_347#_M1017_d N_A_733_66#_M1017_g N_A_1576_99#_M1036_d VPB
+ PHIGHVT L=0.25 W=1 AD=0.23015 AS=0.225 PD=1.51 PS=1.45 NRD=16.0752 NRS=24.6053
+ M=1 R=4 SA=125003 SB=125002 A=0.25 P=2.5 MULT=1
MM1033 A_2095_361# N_A_998_347#_M1033_g N_A_1957_347#_M1017_d VPB PHIGHVT L=0.25
+ W=1 AD=0.1325 AS=0.23015 PD=1.265 PS=1.51 NRD=15.2478 NRS=16.0752 M=1 R=4
+ SA=125003 SB=125001 A=0.25 P=2.5 MULT=1
MM1026 N_VPWR_M1026_d N_A_2148_185#_M1026_g A_2095_361# VPB PHIGHVT L=0.25 W=1
+ AD=0.1775 AS=0.1325 PD=1.355 PS=1.265 NRD=0 NRS=15.2478 M=1 R=4 SA=125004
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1031 N_A_2148_185#_M1031_d N_A_1957_347#_M1031_g N_VPWR_M1026_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.1775 PD=2.57 PS=1.355 NRD=0 NRS=14.7553 M=1 R=4
+ SA=125004 SB=125000 A=0.25 P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_A_2148_185#_M1006_g N_Q_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX38_noxref VNB VPB NWDIODE A=27.3799 P=32.53
*
.include "sky130_fd_sc_lp__sdfxtp_lp.pxi.spice"
*
.ends
*
*
