* File: sky130_fd_sc_lp__a311o_0.pex.spice
* Created: Fri Aug 28 09:57:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311O_0%A_72_312# 1 2 3 12 16 20 21 24 25 27 28 31
+ 33 34 36 41 45 47 48 50 51
r108 50 51 8.96717 $w=4.33e-07 $l=1.85e-07 $layer=LI1_cond $X=3.237 $Y=2.575
+ $X2=3.237 $Y2=2.39
r109 43 45 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.51 $Y=0.74
+ $X2=3.51 $Y2=0.45
r110 42 47 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.2 $Y=0.825 $X2=3.1
+ $Y2=0.825
r111 41 43 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.375 $Y=0.825
+ $X2=3.51 $Y2=0.74
r112 41 42 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.375 $Y=0.825
+ $X2=3.2 $Y2=0.825
r113 37 48 5.27864 $w=1.9e-07 $l=1.02879e-07 $layer=LI1_cond $X=3.11 $Y=2.23
+ $X2=3.1 $Y2=2.132
r114 37 51 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=3.11 $Y=2.23
+ $X2=3.11 $Y2=2.39
r115 36 48 5.27864 $w=1.9e-07 $l=9.7e-08 $layer=LI1_cond $X=3.1 $Y=2.035 $X2=3.1
+ $Y2=2.132
r116 35 47 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.91 $X2=3.1
+ $Y2=0.825
r117 35 36 62.3864 $w=1.98e-07 $l=1.125e-06 $layer=LI1_cond $X=3.1 $Y=0.91
+ $X2=3.1 $Y2=2.035
r118 33 47 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3 $Y=0.825 $X2=3.1
+ $Y2=0.825
r119 33 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3 $Y=0.825
+ $X2=2.725 $Y2=0.825
r120 29 34 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=2.602 $Y=0.74
+ $X2=2.725 $Y2=0.825
r121 29 31 13.6412 $w=2.43e-07 $l=2.9e-07 $layer=LI1_cond $X=2.602 $Y=0.74
+ $X2=2.602 $Y2=0.45
r122 27 48 1.24919 $w=1.95e-07 $l=1e-07 $layer=LI1_cond $X=3 $Y=2.132 $X2=3.1
+ $Y2=2.132
r123 27 28 131.385 $w=1.93e-07 $l=2.31e-06 $layer=LI1_cond $X=3 $Y=2.132
+ $X2=0.69 $Y2=2.132
r124 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.725 $X2=0.525 $Y2=1.725
r125 22 28 6.999 $w=1.95e-07 $l=1.71785e-07 $layer=LI1_cond $X=0.56 $Y=2.035
+ $X2=0.69 $Y2=2.132
r126 22 24 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=0.56 $Y=2.035
+ $X2=0.56 $Y2=1.725
r127 20 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=2.065
+ $X2=0.525 $Y2=1.725
r128 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=2.065
+ $X2=0.525 $Y2=2.23
r129 19 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.56
+ $X2=0.525 $Y2=1.725
r130 16 21 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.615 $Y=2.75
+ $X2=0.615 $Y2=2.23
r131 12 19 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.615 $Y=0.45
+ $X2=0.615 $Y2=1.56
r132 3 50 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.15
+ $Y=2.43 $X2=3.29 $Y2=2.575
r133 2 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.34
+ $Y=0.24 $X2=3.48 $Y2=0.45
r134 1 31 182 $w=1.7e-07 $l=4.99074e-07 $layer=licon1_NDIFF $count=1 $X=2.19
+ $Y=0.24 $X2=2.595 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%A3 3 7 9 10 11 12 13 14 19
c41 19 0 1.01934e-19 $X=1.065 $Y=0.935
c42 3 0 3.97977e-20 $X=1.045 $Y=2.75
r43 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=0.935 $X2=1.065 $Y2=0.935
r44 13 14 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.172 $Y=1.295
+ $X2=1.172 $Y2=1.665
r45 13 20 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=1.172 $Y=1.295
+ $X2=1.172 $Y2=0.935
r46 12 20 0.299336 $w=3.83e-07 $l=1e-08 $layer=LI1_cond $X=1.172 $Y=0.925
+ $X2=1.172 $Y2=0.935
r47 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.065 $Y=1.275
+ $X2=1.065 $Y2=0.935
r48 10 11 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.275
+ $X2=1.065 $Y2=1.44
r49 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=0.77
+ $X2=1.065 $Y2=0.935
r50 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.155 $Y=0.45
+ $X2=1.155 $Y2=0.77
r51 3 11 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=1.045 $Y=2.75
+ $X2=1.045 $Y2=1.44
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%A2 2 5 9 10 11 12 13 14 20 22
r46 20 22 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=0.935
+ $X2=1.62 $Y2=0.77
r47 13 14 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.682 $Y=1.295
+ $X2=1.682 $Y2=1.665
r48 12 13 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.682 $Y=0.925
+ $X2=1.682 $Y2=1.295
r49 12 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.635
+ $Y=0.935 $X2=1.635 $Y2=0.935
r50 11 12 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.682 $Y=0.555
+ $X2=1.682 $Y2=0.925
r51 9 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.575 $Y=0.45
+ $X2=1.575 $Y2=0.77
r52 5 10 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=1.515 $Y=2.75
+ $X2=1.515 $Y2=1.44
r53 2 10 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.62 $Y=1.26 $X2=1.62
+ $Y2=1.44
r54 1 20 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.62 $Y=0.95 $X2=1.62
+ $Y2=0.935
r55 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.62 $Y=0.95 $X2=1.62
+ $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%A1 3 7 11 12 13 14 15 16 22
c47 13 0 9.80436e-20 $X=2.16 $Y=0.555
r48 15 16 16.6906 $w=2.88e-07 $l=4.2e-07 $layer=LI1_cond $X=2.145 $Y=1.245
+ $X2=2.145 $Y2=1.665
r49 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.205
+ $Y=1.245 $X2=2.205 $Y2=1.245
r50 14 15 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=2.145 $Y=0.925
+ $X2=2.145 $Y2=1.245
r51 13 14 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.145 $Y=0.555
+ $X2=2.145 $Y2=0.925
r52 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.205 $Y=1.585
+ $X2=2.205 $Y2=1.245
r53 11 12 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.585
+ $X2=2.205 $Y2=1.75
r54 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.08
+ $X2=2.205 $Y2=1.245
r55 7 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.285 $Y=2.75 $X2=2.285
+ $Y2=1.75
r56 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.115 $Y=0.45
+ $X2=2.115 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%B1 3 7 11 12 13 14 18 19
c46 3 0 1.727e-19 $X=2.715 $Y=2.75
r47 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.745
+ $Y=1.245 $X2=2.745 $Y2=1.245
r48 13 14 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=1.295
+ $X2=2.645 $Y2=1.665
r49 13 19 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=2.645 $Y=1.295
+ $X2=2.645 $Y2=1.245
r50 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.745 $Y=1.585
+ $X2=2.745 $Y2=1.245
r51 11 12 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.585
+ $X2=2.745 $Y2=1.75
r52 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.08
+ $X2=2.745 $Y2=1.245
r53 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.835 $Y=0.45
+ $X2=2.835 $Y2=1.08
r54 3 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.715 $Y=2.75 $X2=2.715
+ $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%C1 3 9 11 12 13 14 15 20
c40 13 0 7.46567e-20 $X=3.6 $Y=1.295
r41 20 22 47.4991 $w=4.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.385 $Y=1.635
+ $X2=3.385 $Y2=1.47
r42 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.455
+ $Y=1.635 $X2=3.455 $Y2=1.635
r43 14 15 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.562 $Y=1.665
+ $X2=3.562 $Y2=2.035
r44 14 21 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=3.562 $Y=1.665
+ $X2=3.562 $Y2=1.635
r45 13 21 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=3.562 $Y=1.295
+ $X2=3.562 $Y2=1.635
r46 11 12 45.7242 $w=4.7e-07 $l=1.5e-07 $layer=POLY_cond $X=3.31 $Y=1.99
+ $X2=3.31 $Y2=2.14
r47 9 22 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.265 $Y=0.45
+ $X2=3.265 $Y2=1.47
r48 5 20 8.28314 $w=4.7e-07 $l=7e-08 $layer=POLY_cond $X=3.385 $Y=1.705
+ $X2=3.385 $Y2=1.635
r49 5 11 33.7242 $w=4.7e-07 $l=2.85e-07 $layer=POLY_cond $X=3.385 $Y=1.705
+ $X2=3.385 $Y2=1.99
r50 3 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.075 $Y=2.75
+ $X2=3.075 $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%X 1 2 10 11 13 14 15 21
r27 15 29 7.45085 $w=4.78e-07 $l=9.5e-08 $layer=LI1_cond $X=0.325 $Y=1.295
+ $X2=0.325 $Y2=1.39
r28 15 19 3.61315 $w=4.78e-07 $l=1.45e-07 $layer=LI1_cond $X=0.325 $Y=1.295
+ $X2=0.325 $Y2=1.15
r29 14 19 5.60662 $w=4.78e-07 $l=2.25e-07 $layer=LI1_cond $X=0.325 $Y=0.925
+ $X2=0.325 $Y2=1.15
r30 13 14 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.325 $Y=0.555
+ $X2=0.325 $Y2=0.925
r31 13 21 2.61642 $w=4.78e-07 $l=1.05e-07 $layer=LI1_cond $X=0.325 $Y=0.555
+ $X2=0.325 $Y2=0.45
r32 11 29 64.6442 $w=1.73e-07 $l=1.02e-06 $layer=LI1_cond $X=0.172 $Y=2.41
+ $X2=0.172 $Y2=1.39
r33 10 11 9.19513 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.325 $Y=2.575
+ $X2=0.325 $Y2=2.41
r34 2 10 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.255
+ $Y=2.43 $X2=0.4 $Y2=2.575
r35 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.24 $X2=0.4 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%VPWR 1 2 9 11 13 14 15 23 24 27
r42 30 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 27 30 9.5912 $w=5.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.9 $Y=2.905 $X2=1.9
+ $Y2=3.33
r45 24 33 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 21 30 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=1.9 $Y2=3.33
r48 21 23 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 19 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 15 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 15 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 13 18 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 13 14 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.85 $Y2=3.33
r55 12 14 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.85 $Y2=3.33
r56 11 30 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=1.9 $Y2=3.33
r57 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=0.965 $Y2=3.33
r58 7 14 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=3.33
r59 7 9 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=0.85 $Y=3.245 $X2=0.85
+ $Y2=2.575
r60 2 27 300 $w=1.7e-07 $l=6.77052e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=2.43 $X2=2.07 $Y2=2.905
r61 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=2.43 $X2=0.83 $Y2=2.575
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%A_224_486# 1 2 9 11 12 15
c29 9 0 3.97977e-20 $X=1.3 $Y=2.575
r30 13 15 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.5 $Y=2.57 $X2=2.5
+ $Y2=2.575
r31 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=2.485
+ $X2=2.5 $Y2=2.57
r32 11 12 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.335 $Y=2.485
+ $X2=1.465 $Y2=2.485
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.3 $Y=2.57
+ $X2=1.465 $Y2=2.485
r34 7 9 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.3 $Y=2.57 $X2=1.3
+ $Y2=2.575
r35 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=2.43 $X2=2.5 $Y2=2.575
r36 1 9 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=1.12
+ $Y=2.43 $X2=1.3 $Y2=2.575
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_0%VGND 1 2 9 13 16 17 18 24 33 34 37
c51 24 0 1.01934e-19 $X=2.895 $Y=0
r52 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 34 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r54 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 31 37 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.05
+ $Y2=0
r56 31 33 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.6
+ $Y2=0
r57 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r58 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r59 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r60 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 24 37 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=3.05
+ $Y2=0
r62 24 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=2.64
+ $Y2=0
r63 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r64 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 18 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r66 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r67 16 21 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.72
+ $Y2=0
r68 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=0 $X2=0.9
+ $Y2=0
r69 15 26 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.2
+ $Y2=0
r70 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.9
+ $Y2=0
r71 11 37 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0
r72 11 13 11.8962 $w=3.08e-07 $l=3.2e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0.405
r73 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0
r74 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.9 $Y=0.085 $X2=0.9
+ $Y2=0.435
r75 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.91
+ $Y=0.24 $X2=3.05 $Y2=0.405
r76 1 9 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.24 $X2=0.9 $Y2=0.435
.ends

