* File: sky130_fd_sc_lp__xor2_1.spice
* Created: Wed Sep  2 10:41:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor2_1.pex.spice"
.subckt sky130_fd_sc_lp__xor2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1008 N_A_42_367#_M1008_d N_B_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_42_367#_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1002 A_297_69# N_A_M1002_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.1176 PD=1.08 PS=1.12 NRD=9.276 NRS=0 M=1 R=5.6 SA=75001.1 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1003 N_X_M1003_d N_B_M1003_g A_297_69# VNB NSHORT L=0.15 W=0.84 AD=0.2436
+ AS=0.1008 PD=1.42 PS=1.08 NRD=27.132 NRS=9.276 M=1 R=5.6 SA=75001.4 SB=75001.2
+ A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A_42_367#_M1000_g N_X_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.4788 AS=0.2436 PD=2.82 PS=1.42 NRD=43.56 NRS=15.708 M=1 R=5.6 SA=75002.2
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1001 A_125_367# N_B_M1001_g N_A_42_367#_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3339 PD=1.5 PS=3.05 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_125_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.1512 PD=1.56 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6 SB=75001.2
+ A=0.189 P=2.82 MULT=1
MM1007 N_A_293_367#_M1007_d N_A_M1007_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.189 PD=1.54 PS=1.56 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75001
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_293_367#_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4786 AS=0.1764 PD=3.44 PS=1.54 NRD=15.6221 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.3 A=0.189 P=2.82 MULT=1
MM1005 N_A_293_367#_M1005_d N_A_42_367#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3591 PD=3.05 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__xor2_1.pxi.spice"
*
.ends
*
*
