* File: sky130_fd_sc_lp__mux4_m.pxi.spice
* Created: Fri Aug 28 10:46:37 2020
* 
x_PM_SKY130_FD_SC_LP__MUX4_M%A2 N_A2_M1001_g N_A2_M1024_g N_A2_c_180_n
+ N_A2_c_181_n A2 A2 A2 A2 N_A2_c_178_n PM_SKY130_FD_SC_LP__MUX4_M%A2
x_PM_SKY130_FD_SC_LP__MUX4_M%A_59_463# N_A_59_463#_M1014_s N_A_59_463#_M1023_s
+ N_A_59_463#_M1020_g N_A_59_463#_M1013_g N_A_59_463#_M1004_g
+ N_A_59_463#_M1016_g N_A_59_463#_c_217_n N_A_59_463#_c_218_n
+ N_A_59_463#_c_236_n N_A_59_463#_c_219_n N_A_59_463#_c_220_n
+ N_A_59_463#_c_221_n N_A_59_463#_c_222_n N_A_59_463#_c_223_n
+ N_A_59_463#_c_224_n N_A_59_463#_c_225_n N_A_59_463#_c_226_n
+ N_A_59_463#_c_227_n N_A_59_463#_c_228_n N_A_59_463#_c_229_n
+ N_A_59_463#_c_230_n N_A_59_463#_c_231_n N_A_59_463#_c_232_n
+ PM_SKY130_FD_SC_LP__MUX4_M%A_59_463#
x_PM_SKY130_FD_SC_LP__MUX4_M%A3 N_A3_M1007_g N_A3_M1003_g N_A3_c_361_n
+ N_A3_c_366_n A3 N_A3_c_363_n PM_SKY130_FD_SC_LP__MUX4_M%A3
x_PM_SKY130_FD_SC_LP__MUX4_M%A1 N_A1_M1022_g N_A1_M1011_g N_A1_c_406_n
+ N_A1_c_410_n A1 N_A1_c_407_n N_A1_c_420_n PM_SKY130_FD_SC_LP__MUX4_M%A1
x_PM_SKY130_FD_SC_LP__MUX4_M%S0 N_S0_M1023_g N_S0_M1014_g N_S0_c_449_n
+ N_S0_M1000_g N_S0_c_463_n N_S0_c_464_n N_S0_M1006_g N_S0_c_451_n N_S0_M1015_g
+ N_S0_c_453_n N_S0_M1017_g N_S0_c_466_n N_S0_c_454_n N_S0_c_455_n N_S0_c_456_n
+ N_S0_c_457_n N_S0_c_468_n N_S0_c_458_n S0 N_S0_c_459_n N_S0_c_460_n
+ PM_SKY130_FD_SC_LP__MUX4_M%S0
x_PM_SKY130_FD_SC_LP__MUX4_M%A0 N_A0_c_582_n N_A0_M1009_g N_A0_M1019_g A0
+ N_A0_c_585_n PM_SKY130_FD_SC_LP__MUX4_M%A0
x_PM_SKY130_FD_SC_LP__MUX4_M%A_1118_37# N_A_1118_37#_M1025_s
+ N_A_1118_37#_M1010_s N_A_1118_37#_M1018_g N_A_1118_37#_c_619_n
+ N_A_1118_37#_M1005_g N_A_1118_37#_c_616_n N_A_1118_37#_c_617_n
+ N_A_1118_37#_c_621_n N_A_1118_37#_c_622_n N_A_1118_37#_c_623_n
+ N_A_1118_37#_c_643_p N_A_1118_37#_c_624_n
+ PM_SKY130_FD_SC_LP__MUX4_M%A_1118_37#
x_PM_SKY130_FD_SC_LP__MUX4_M%S1 N_S1_M1012_g N_S1_c_694_n N_S1_c_695_n
+ N_S1_c_685_n N_S1_M1021_g N_S1_c_686_n N_S1_c_687_n N_S1_c_696_n N_S1_c_688_n
+ N_S1_c_689_n N_S1_M1025_g N_S1_c_698_n N_S1_M1010_g N_S1_c_699_n N_S1_c_690_n
+ N_S1_c_691_n S1 N_S1_c_692_n PM_SKY130_FD_SC_LP__MUX4_M%S1
x_PM_SKY130_FD_SC_LP__MUX4_M%A_1184_171# N_A_1184_171#_M1018_d
+ N_A_1184_171#_M1012_d N_A_1184_171#_c_769_n N_A_1184_171#_M1008_g
+ N_A_1184_171#_M1002_g N_A_1184_171#_c_771_n N_A_1184_171#_c_778_n
+ N_A_1184_171#_c_772_n N_A_1184_171#_c_780_n N_A_1184_171#_c_773_n
+ N_A_1184_171#_c_774_n N_A_1184_171#_c_775_n N_A_1184_171#_c_782_n
+ PM_SKY130_FD_SC_LP__MUX4_M%A_1184_171#
x_PM_SKY130_FD_SC_LP__MUX4_M%VPWR N_VPWR_M1023_d N_VPWR_M1007_d N_VPWR_M1019_d
+ N_VPWR_M1010_d N_VPWR_c_831_n N_VPWR_c_832_n N_VPWR_c_833_n N_VPWR_c_834_n
+ N_VPWR_c_835_n N_VPWR_c_836_n N_VPWR_c_837_n N_VPWR_c_838_n VPWR
+ N_VPWR_c_839_n N_VPWR_c_840_n N_VPWR_c_841_n N_VPWR_c_830_n N_VPWR_c_843_n
+ N_VPWR_c_844_n PM_SKY130_FD_SC_LP__MUX4_M%VPWR
x_PM_SKY130_FD_SC_LP__MUX4_M%A_345_126# N_A_345_126#_M1020_d
+ N_A_345_126#_M1021_d N_A_345_126#_M1000_d N_A_345_126#_M1005_d
+ N_A_345_126#_c_974_n N_A_345_126#_c_914_n N_A_345_126#_c_921_n
+ N_A_345_126#_c_922_n N_A_345_126#_c_951_n N_A_345_126#_c_923_n
+ N_A_345_126#_c_924_n N_A_345_126#_c_925_n N_A_345_126#_c_926_n
+ N_A_345_126#_c_927_n N_A_345_126#_c_928_n N_A_345_126#_c_929_n
+ N_A_345_126#_c_930_n N_A_345_126#_c_915_n N_A_345_126#_c_916_n
+ N_A_345_126#_c_917_n N_A_345_126#_c_932_n N_A_345_126#_c_918_n
+ N_A_345_126#_c_933_n N_A_345_126#_c_919_n N_A_345_126#_c_934_n
+ PM_SKY130_FD_SC_LP__MUX4_M%A_345_126#
x_PM_SKY130_FD_SC_LP__MUX4_M%A_688_126# N_A_688_126#_M1015_d
+ N_A_688_126#_M1018_s N_A_688_126#_M1004_d N_A_688_126#_M1012_s
+ N_A_688_126#_c_1080_n N_A_688_126#_c_1083_n N_A_688_126#_c_1071_n
+ N_A_688_126#_c_1074_n N_A_688_126#_c_1075_n N_A_688_126#_c_1072_n
+ N_A_688_126#_c_1077_n N_A_688_126#_c_1078_n N_A_688_126#_c_1079_n
+ PM_SKY130_FD_SC_LP__MUX4_M%A_688_126#
x_PM_SKY130_FD_SC_LP__MUX4_M%X N_X_M1008_d N_X_M1002_d X X X X X X N_X_c_1132_n
+ PM_SKY130_FD_SC_LP__MUX4_M%X
x_PM_SKY130_FD_SC_LP__MUX4_M%VGND N_VGND_M1014_d N_VGND_M1003_d N_VGND_M1009_d
+ N_VGND_M1025_d N_VGND_c_1145_n N_VGND_c_1146_n N_VGND_c_1147_n N_VGND_c_1148_n
+ N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n N_VGND_c_1152_n VGND
+ N_VGND_c_1153_n N_VGND_c_1154_n N_VGND_c_1155_n N_VGND_c_1156_n
+ N_VGND_c_1157_n N_VGND_c_1158_n PM_SKY130_FD_SC_LP__MUX4_M%VGND
cc_1 VNB N_A2_M1001_g 0.0322937f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.84
cc_2 VNB A2 9.47981e-19 $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_3 VNB N_A2_c_178_n 0.0169634f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.65
cc_4 VNB N_A_59_463#_M1016_g 0.0391292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_59_463#_c_217_n 0.0133923f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.65
cc_6 VNB N_A_59_463#_c_218_n 0.0232721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_59_463#_c_219_n 0.0172407f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.775
cc_8 VNB N_A_59_463#_c_220_n 0.0249949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_59_463#_c_221_n 0.00281366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_59_463#_c_222_n 0.00292383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_59_463#_c_223_n 0.0180474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_59_463#_c_224_n 0.0167603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_59_463#_c_225_n 0.00276201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_59_463#_c_226_n 0.00235244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_59_463#_c_227_n 0.0329468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_59_463#_c_228_n 0.002243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_59_463#_c_229_n 0.00485122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_59_463#_c_230_n 0.0219604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_59_463#_c_231_n 0.00420897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_59_463#_c_232_n 0.0167535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_M1003_g 0.0261197f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=2.525
cc_22 VNB N_A3_c_361_n 0.00637713f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.99
cc_23 VNB A3 0.00278471f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_24 VNB N_A3_c_363_n 0.0162224f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.69
cc_25 VNB N_A1_M1022_g 0.0279339f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.84
cc_26 VNB N_A1_c_406_n 0.00675672f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.99
cc_27 VNB N_A1_c_407_n 0.0173763f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.69
cc_28 VNB N_S0_M1023_g 0.020925f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.84
cc_29 VNB N_S0_M1014_g 0.0144355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_S0_c_449_n 0.0910467f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.65
cc_31 VNB N_S0_M1006_g 0.0368778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_S0_c_451_n 0.0742047f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.65
cc_33 VNB N_S0_M1015_g 0.0380117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_S0_c_453_n 0.119705f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.035
cc_35 VNB N_S0_c_454_n 0.0950502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_S0_c_455_n 0.0200817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_S0_c_456_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_S0_c_457_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_S0_c_458_n 8.79809e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_S0_c_459_n 0.0645807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_S0_c_460_n 0.0228343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A0_c_582_n 0.0173612f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.485
cc_43 VNB N_A0_M1019_g 0.010413f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=2.525
cc_44 VNB A0 0.00707277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A0_c_585_n 0.0464775f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.99
cc_46 VNB N_A_1118_37#_M1018_g 0.0511752f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.485
cc_47 VNB N_A_1118_37#_c_616_n 0.0288304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1118_37#_c_617_n 0.0480199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_S1_c_685_n 0.017914f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=2.525
cc_50 VNB N_S1_c_686_n 0.0245938f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.485
cc_51 VNB N_S1_c_687_n 0.00817669f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.99
cc_52 VNB N_S1_c_688_n 0.00413229f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.32
cc_53 VNB N_S1_c_689_n 0.0204383f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.69
cc_54 VNB N_S1_c_690_n 0.032601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_S1_c_691_n 0.0124659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_S1_c_692_n 0.0356649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1184_171#_c_769_n 0.0214981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1184_171#_M1008_g 0.0454328f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.99
cc_59 VNB N_A_1184_171#_c_771_n 0.00569649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1184_171#_c_772_n 0.0139017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1184_171#_c_773_n 0.00363798f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.405
cc_62 VNB N_A_1184_171#_c_774_n 0.0244091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1184_171#_c_775_n 0.00128461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VPWR_c_830_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_345_126#_c_914_n 0.00843817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_345_126#_c_915_n 0.00389725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_345_126#_c_916_n 0.0148069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_345_126#_c_917_n 0.00363776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_345_126#_c_918_n 0.00134984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_345_126#_c_919_n 0.00171982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_688_126#_c_1071_n 0.0120118f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.65
cc_72 VNB N_A_688_126#_c_1072_n 0.00901363f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.405
cc_73 VNB N_X_c_1132_n 0.050724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1145_n 0.00985612f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.32
cc_75 VNB N_VGND_c_1146_n 0.00846146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1147_n 0.0182243f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.65
cc_77 VNB N_VGND_c_1148_n 0.00482866f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.035
cc_78 VNB N_VGND_c_1149_n 0.0363432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1150_n 0.00256535f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.775
cc_80 VNB N_VGND_c_1151_n 0.039093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1152_n 0.00283539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1153_n 0.0243474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1154_n 0.0772085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1155_n 0.0191183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1156_n 0.424799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1157_n 0.00445561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1158_n 0.00362723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VPB N_A2_M1024_g 0.020087f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=2.525
cc_89 VPB N_A2_c_180_n 0.0265814f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.99
cc_90 VPB N_A2_c_181_n 0.0216239f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.155
cc_91 VPB A2 0.00363855f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_92 VPB N_A_59_463#_M1013_g 0.0341777f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.155
cc_93 VPB N_A_59_463#_M1004_g 0.0320414f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.69
cc_94 VPB N_A_59_463#_c_218_n 0.00168511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_59_463#_c_236_n 0.0309867f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.035
cc_96 VPB N_A_59_463#_c_219_n 0.0343268f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_97 VPB N_A_59_463#_c_222_n 0.00757855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_59_463#_c_229_n 0.0014395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_59_463#_c_232_n 0.0274279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A3_M1007_g 0.0229483f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=0.84
cc_101 VPB N_A3_c_361_n 0.01346f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.99
cc_102 VPB N_A3_c_366_n 0.0147573f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.155
cc_103 VPB A3 0.0043984f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_104 VPB N_A1_M1011_g 0.0221858f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=2.525
cc_105 VPB N_A1_c_406_n 0.0163128f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.99
cc_106 VPB N_A1_c_410_n 0.0158635f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.155
cc_107 VPB N_S0_M1023_g 0.0551188f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=0.84
cc_108 VPB N_S0_M1000_g 0.036354f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_109 VPB N_S0_c_463_n 0.157622f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.32
cc_110 VPB N_S0_c_464_n 0.0126165f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.69
cc_111 VPB N_S0_M1017_g 0.0336821f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_112 VPB N_S0_c_466_n 0.0731925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_S0_c_454_n 0.0956588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_S0_c_468_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A0_M1019_g 0.0457276f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=2.525
cc_116 VPB N_A_1118_37#_M1018_g 0.00915057f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.485
cc_117 VPB N_A_1118_37#_c_619_n 0.00926484f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.155
cc_118 VPB N_A_1118_37#_M1005_g 0.0197323f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.32
cc_119 VPB N_A_1118_37#_c_621_n 0.00742661f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.65
cc_120 VPB N_A_1118_37#_c_622_n 0.0472393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_1118_37#_c_623_n 0.00983104f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.405
cc_122 VPB N_A_1118_37#_c_624_n 0.022752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_S1_M1012_g 0.0376324f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=0.84
cc_124 VPB N_S1_c_694_n 0.0608832f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=2.155
cc_125 VPB N_S1_c_695_n 0.012806f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=2.525
cc_126 VPB N_S1_c_696_n 0.0335241f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_127 VPB N_S1_c_688_n 0.0377153f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.32
cc_128 VPB N_S1_c_698_n 0.0172234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_S1_c_699_n 0.0367033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_1184_171#_c_769_n 5.38414e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_1184_171#_M1002_g 0.0610398f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.32
cc_132 VPB N_A_1184_171#_c_778_n 0.0109819f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.65
cc_133 VPB N_A_1184_171#_c_772_n 0.0108815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_1184_171#_c_780_n 0.00666727f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.035
cc_135 VPB N_A_1184_171#_c_775_n 3.01005e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_1184_171#_c_782_n 0.0252649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_831_n 0.0205482f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.32
cc_138 VPB N_VPWR_c_832_n 0.0163483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_833_n 0.00940455f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.65
cc_140 VPB N_VPWR_c_834_n 0.00606944f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.035
cc_141 VPB N_VPWR_c_835_n 0.0250453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_836_n 0.00362871f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_143 VPB N_VPWR_c_837_n 0.0439875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_838_n 0.00223798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_839_n 0.0465286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_840_n 0.0678343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_841_n 0.0192421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_830_n 0.102077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_843_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_844_n 0.00401309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_345_126#_c_914_n 0.00413972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_345_126#_c_921_n 0.0162487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_345_126#_c_922_n 0.00413217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_345_126#_c_923_n 0.024325f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.65
cc_155 VPB N_A_345_126#_c_924_n 0.00239194f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.65
cc_156 VPB N_A_345_126#_c_925_n 0.00119894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_345_126#_c_926_n 0.018848f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.035
cc_158 VPB N_A_345_126#_c_927_n 0.00142255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_345_126#_c_928_n 0.00485606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_345_126#_c_929_n 0.0208825f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.775
cc_161 VPB N_A_345_126#_c_930_n 7.35373e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_345_126#_c_915_n 0.00742247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_345_126#_c_932_n 0.0110298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_345_126#_c_933_n 0.00122223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_345_126#_c_934_n 0.00124581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_688_126#_c_1071_n 0.00150463f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.65
cc_167 VPB N_A_688_126#_c_1074_n 0.00690969f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.65
cc_168 VPB N_A_688_126#_c_1075_n 0.0389562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_688_126#_c_1072_n 0.0016495f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=2.405
cc_170 VPB N_A_688_126#_c_1077_n 0.00942742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_688_126#_c_1078_n 0.00215798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_688_126#_c_1079_n 0.00312145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_X_c_1132_n 0.0505796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 N_A2_c_180_n N_A_59_463#_M1013_g 0.00691667f $X=1.2 $Y=1.99 $X2=0 $Y2=0
cc_175 N_A2_M1001_g N_A_59_463#_c_217_n 0.0267687f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_176 N_A2_c_180_n N_A_59_463#_c_218_n 0.0267687f $X=1.2 $Y=1.99 $X2=0 $Y2=0
cc_177 A2 N_A_59_463#_c_218_n 3.49949e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_178 A2 N_A_59_463#_c_219_n 0.0255583f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A2_M1001_g N_A_59_463#_c_220_n 0.0173593f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_180 A2 N_A_59_463#_c_220_n 0.0125942f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A2_c_178_n N_A_59_463#_c_220_n 0.00397544f $X=1.2 $Y=1.65 $X2=0 $Y2=0
cc_182 N_A2_M1001_g N_A_59_463#_c_221_n 0.00364681f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_183 N_A2_M1001_g N_A_59_463#_c_222_n 0.0063734f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_184 A2 N_A_59_463#_c_222_n 0.0203113f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A2_c_178_n N_A_59_463#_c_223_n 0.0267687f $X=1.2 $Y=1.65 $X2=0 $Y2=0
cc_186 N_A2_M1001_g N_A_59_463#_c_230_n 0.0010586f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_187 N_A2_M1001_g N_S0_M1023_g 0.00439528f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_188 N_A2_M1024_g N_S0_M1023_g 0.00968493f $X=1.29 $Y=2.525 $X2=0 $Y2=0
cc_189 A2 N_S0_M1023_g 0.00490855f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_190 N_A2_c_178_n N_S0_M1023_g 0.0242365f $X=1.2 $Y=1.65 $X2=0 $Y2=0
cc_191 N_A2_M1001_g N_S0_c_449_n 0.00908269f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_192 N_A2_M1024_g N_S0_M1000_g 0.0395871f $X=1.29 $Y=2.525 $X2=0 $Y2=0
cc_193 A2 N_S0_M1000_g 0.00265441f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A2_M1001_g N_S0_c_459_n 0.016566f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_195 A2 N_VPWR_M1023_d 0.00463432f $X=1.115 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_196 N_A2_M1024_g N_VPWR_c_831_n 0.00141151f $X=1.29 $Y=2.525 $X2=0 $Y2=0
cc_197 A2 N_VPWR_c_831_n 0.0308777f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A2_M1024_g N_VPWR_c_839_n 0.00380937f $X=1.29 $Y=2.525 $X2=0 $Y2=0
cc_199 A2 N_VPWR_c_839_n 0.00485955f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A2_M1024_g N_VPWR_c_830_n 0.00477801f $X=1.29 $Y=2.525 $X2=0 $Y2=0
cc_201 A2 N_VPWR_c_830_n 0.00566862f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_202 N_A2_c_180_n N_A_345_126#_c_914_n 0.00189266f $X=1.2 $Y=1.99 $X2=0 $Y2=0
cc_203 N_A2_M1024_g N_A_345_126#_c_922_n 3.54487e-19 $X=1.29 $Y=2.525 $X2=0
+ $Y2=0
cc_204 A2 N_A_345_126#_c_922_n 0.00560127f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A2_M1001_g N_VGND_c_1145_n 0.00159777f $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_206 N_A2_M1001_g N_VGND_c_1156_n 9.43998e-19 $X=1.29 $Y=0.84 $X2=0 $Y2=0
cc_207 N_A_59_463#_c_223_n N_A3_M1003_g 0.00284068f $X=1.74 $Y=1.325 $X2=0 $Y2=0
cc_208 N_A_59_463#_c_226_n N_A3_M1003_g 0.011874f $X=2.44 $Y=1.1 $X2=0 $Y2=0
cc_209 N_A_59_463#_c_227_n N_A3_M1003_g 0.0093486f $X=3.525 $Y=1.185 $X2=0 $Y2=0
cc_210 N_A_59_463#_c_228_n N_A3_M1003_g 0.00302571f $X=2.525 $Y=1.185 $X2=0
+ $Y2=0
cc_211 N_A_59_463#_c_236_n N_A3_c_361_n 0.0367909f $X=2.08 $Y=1.755 $X2=0 $Y2=0
cc_212 N_A_59_463#_M1013_g N_A3_c_366_n 0.0367909f $X=2.08 $Y=2.525 $X2=0 $Y2=0
cc_213 N_A_59_463#_c_236_n A3 3.61298e-19 $X=2.08 $Y=1.755 $X2=0 $Y2=0
cc_214 N_A_59_463#_c_227_n A3 0.0134794f $X=3.525 $Y=1.185 $X2=0 $Y2=0
cc_215 N_A_59_463#_c_228_n A3 0.0120394f $X=2.525 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A_59_463#_c_218_n N_A3_c_363_n 0.00582674f $X=1.74 $Y=1.68 $X2=0 $Y2=0
cc_217 N_A_59_463#_c_227_n N_A3_c_363_n 0.001954f $X=3.525 $Y=1.185 $X2=0 $Y2=0
cc_218 N_A_59_463#_c_228_n N_A3_c_363_n 0.00324021f $X=2.525 $Y=1.185 $X2=0
+ $Y2=0
cc_219 N_A_59_463#_M1016_g N_A1_M1022_g 0.00225459f $X=3.795 $Y=0.84 $X2=0 $Y2=0
cc_220 N_A_59_463#_c_226_n N_A1_M1022_g 9.7207e-19 $X=2.44 $Y=1.1 $X2=0 $Y2=0
cc_221 N_A_59_463#_c_227_n N_A1_M1022_g 0.0155263f $X=3.525 $Y=1.185 $X2=0 $Y2=0
cc_222 N_A_59_463#_c_229_n N_A1_M1022_g 0.00203691f $X=3.61 $Y=1.715 $X2=0 $Y2=0
cc_223 N_A_59_463#_M1004_g N_A1_c_410_n 0.0402766f $X=3.52 $Y=2.525 $X2=0 $Y2=0
cc_224 N_A_59_463#_M1016_g N_A1_c_407_n 0.00272934f $X=3.795 $Y=0.84 $X2=0 $Y2=0
cc_225 N_A_59_463#_c_227_n N_A1_c_407_n 0.0051156f $X=3.525 $Y=1.185 $X2=0 $Y2=0
cc_226 N_A_59_463#_c_229_n N_A1_c_407_n 0.00329104f $X=3.61 $Y=1.715 $X2=0 $Y2=0
cc_227 N_A_59_463#_c_232_n N_A1_c_407_n 0.0402766f $X=3.795 $Y=1.715 $X2=0 $Y2=0
cc_228 N_A_59_463#_c_227_n N_A1_c_420_n 0.0220798f $X=3.525 $Y=1.185 $X2=0 $Y2=0
cc_229 N_A_59_463#_c_229_n N_A1_c_420_n 0.0193882f $X=3.61 $Y=1.715 $X2=0 $Y2=0
cc_230 N_A_59_463#_c_232_n N_A1_c_420_n 0.00167399f $X=3.795 $Y=1.715 $X2=0
+ $Y2=0
cc_231 N_A_59_463#_c_220_n N_S0_M1014_g 0.00621783f $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_232 N_A_59_463#_c_221_n N_S0_M1014_g 5.42675e-19 $X=1.605 $Y=1.135 $X2=0
+ $Y2=0
cc_233 N_A_59_463#_c_230_n N_S0_M1014_g 0.00881826f $X=0.535 $Y=0.905 $X2=0
+ $Y2=0
cc_234 N_A_59_463#_c_217_n N_S0_c_449_n 0.00739793f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A_59_463#_c_224_n N_S0_c_449_n 0.0072643f $X=2.355 $Y=0.36 $X2=0 $Y2=0
cc_236 N_A_59_463#_c_225_n N_S0_c_449_n 0.00235392f $X=1.69 $Y=0.36 $X2=0 $Y2=0
cc_237 N_A_59_463#_M1013_g N_S0_M1000_g 0.0158604f $X=2.08 $Y=2.525 $X2=0 $Y2=0
cc_238 N_A_59_463#_c_236_n N_S0_M1000_g 0.00520779f $X=2.08 $Y=1.755 $X2=0 $Y2=0
cc_239 N_A_59_463#_c_222_n N_S0_M1000_g 0.00107117f $X=1.74 $Y=1.325 $X2=0 $Y2=0
cc_240 N_A_59_463#_M1013_g N_S0_c_463_n 0.0104164f $X=2.08 $Y=2.525 $X2=0 $Y2=0
cc_241 N_A_59_463#_M1004_g N_S0_c_463_n 0.00889704f $X=3.52 $Y=2.525 $X2=0 $Y2=0
cc_242 N_A_59_463#_c_217_n N_S0_M1006_g 0.0121203f $X=1.74 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_59_463#_c_236_n N_S0_M1006_g 7.81193e-19 $X=2.08 $Y=1.755 $X2=0 $Y2=0
cc_244 N_A_59_463#_c_221_n N_S0_M1006_g 0.00169334f $X=1.605 $Y=1.135 $X2=0
+ $Y2=0
cc_245 N_A_59_463#_c_223_n N_S0_M1006_g 0.00123393f $X=1.74 $Y=1.325 $X2=0 $Y2=0
cc_246 N_A_59_463#_c_224_n N_S0_M1006_g 0.0157725f $X=2.355 $Y=0.36 $X2=0 $Y2=0
cc_247 N_A_59_463#_c_226_n N_S0_M1006_g 0.00559332f $X=2.44 $Y=1.1 $X2=0 $Y2=0
cc_248 N_A_59_463#_c_228_n N_S0_M1006_g 5.44813e-19 $X=2.525 $Y=1.185 $X2=0
+ $Y2=0
cc_249 N_A_59_463#_c_224_n N_S0_c_451_n 0.00339656f $X=2.355 $Y=0.36 $X2=0 $Y2=0
cc_250 N_A_59_463#_M1016_g N_S0_M1015_g 0.0139271f $X=3.795 $Y=0.84 $X2=0 $Y2=0
cc_251 N_A_59_463#_c_227_n N_S0_M1015_g 0.0108636f $X=3.525 $Y=1.185 $X2=0 $Y2=0
cc_252 N_A_59_463#_M1016_g N_S0_c_453_n 0.00846129f $X=3.795 $Y=0.84 $X2=0 $Y2=0
cc_253 N_A_59_463#_M1004_g N_S0_M1017_g 0.0150738f $X=3.52 $Y=2.525 $X2=0 $Y2=0
cc_254 N_A_59_463#_c_219_n N_S0_c_455_n 0.030809f $X=0.42 $Y=2.46 $X2=0 $Y2=0
cc_255 N_A_59_463#_c_220_n N_S0_c_455_n 0.00897463f $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_256 N_A_59_463#_c_230_n N_S0_c_455_n 0.0140127f $X=0.535 $Y=0.905 $X2=0 $Y2=0
cc_257 N_A_59_463#_c_230_n N_S0_c_458_n 0.0115032f $X=0.535 $Y=0.905 $X2=0 $Y2=0
cc_258 N_A_59_463#_c_230_n N_S0_c_459_n 0.00601911f $X=0.535 $Y=0.905 $X2=0
+ $Y2=0
cc_259 N_A_59_463#_c_230_n N_S0_c_460_n 6.66761e-19 $X=0.535 $Y=0.905 $X2=0
+ $Y2=0
cc_260 N_A_59_463#_M1016_g N_A0_c_582_n 0.04615f $X=3.795 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_261 N_A_59_463#_M1004_g N_A0_M1019_g 0.00328171f $X=3.52 $Y=2.525 $X2=0 $Y2=0
cc_262 N_A_59_463#_c_232_n N_A0_M1019_g 0.00760707f $X=3.795 $Y=1.715 $X2=0
+ $Y2=0
cc_263 N_A_59_463#_M1016_g N_A0_c_585_n 0.00760707f $X=3.795 $Y=0.84 $X2=0 $Y2=0
cc_264 N_A_59_463#_M1013_g N_VPWR_c_832_n 0.00146534f $X=2.08 $Y=2.525 $X2=0
+ $Y2=0
cc_265 N_A_59_463#_c_219_n N_VPWR_c_835_n 0.00328868f $X=0.42 $Y=2.46 $X2=0
+ $Y2=0
cc_266 N_A_59_463#_M1013_g N_VPWR_c_830_n 9.39239e-19 $X=2.08 $Y=2.525 $X2=0
+ $Y2=0
cc_267 N_A_59_463#_c_219_n N_VPWR_c_830_n 0.00599347f $X=0.42 $Y=2.46 $X2=0
+ $Y2=0
cc_268 N_A_59_463#_M1013_g N_A_345_126#_c_914_n 0.0118752f $X=2.08 $Y=2.525
+ $X2=0 $Y2=0
cc_269 N_A_59_463#_c_217_n N_A_345_126#_c_914_n 0.00128086f $X=1.74 $Y=1.16
+ $X2=0 $Y2=0
cc_270 N_A_59_463#_c_236_n N_A_345_126#_c_914_n 0.00788309f $X=2.08 $Y=1.755
+ $X2=0 $Y2=0
cc_271 N_A_59_463#_c_221_n N_A_345_126#_c_914_n 0.00798055f $X=1.605 $Y=1.135
+ $X2=0 $Y2=0
cc_272 N_A_59_463#_c_222_n N_A_345_126#_c_914_n 0.0368926f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_273 N_A_59_463#_c_223_n N_A_345_126#_c_914_n 0.00522691f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_274 N_A_59_463#_c_226_n N_A_345_126#_c_914_n 0.00977092f $X=2.44 $Y=1.1 $X2=0
+ $Y2=0
cc_275 N_A_59_463#_c_228_n N_A_345_126#_c_914_n 0.0134815f $X=2.525 $Y=1.185
+ $X2=0 $Y2=0
cc_276 N_A_59_463#_c_231_n N_A_345_126#_c_914_n 0.0131207f $X=1.672 $Y=1.22
+ $X2=0 $Y2=0
cc_277 N_A_59_463#_M1004_g N_A_345_126#_c_921_n 9.70651e-19 $X=3.52 $Y=2.525
+ $X2=0 $Y2=0
cc_278 N_A_59_463#_M1013_g N_A_345_126#_c_922_n 0.0119489f $X=2.08 $Y=2.525
+ $X2=0 $Y2=0
cc_279 N_A_59_463#_c_236_n N_A_345_126#_c_922_n 0.00599027f $X=2.08 $Y=1.755
+ $X2=0 $Y2=0
cc_280 N_A_59_463#_c_222_n N_A_345_126#_c_922_n 0.00300858f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_281 N_A_59_463#_M1004_g N_A_345_126#_c_951_n 0.00174348f $X=3.52 $Y=2.525
+ $X2=0 $Y2=0
cc_282 N_A_59_463#_M1004_g N_A_345_126#_c_923_n 0.0104347f $X=3.52 $Y=2.525
+ $X2=0 $Y2=0
cc_283 N_A_59_463#_c_217_n N_A_345_126#_c_919_n 0.00245f $X=1.74 $Y=1.16 $X2=0
+ $Y2=0
cc_284 N_A_59_463#_c_221_n N_A_345_126#_c_919_n 0.0231944f $X=1.605 $Y=1.135
+ $X2=0 $Y2=0
cc_285 N_A_59_463#_c_223_n N_A_345_126#_c_919_n 0.00148206f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_286 N_A_59_463#_c_224_n N_A_345_126#_c_919_n 0.0213027f $X=2.355 $Y=0.36
+ $X2=0 $Y2=0
cc_287 N_A_59_463#_c_226_n N_A_345_126#_c_919_n 0.0231466f $X=2.44 $Y=1.1 $X2=0
+ $Y2=0
cc_288 N_A_59_463#_M1016_g N_A_688_126#_c_1080_n 0.0136398f $X=3.795 $Y=0.84
+ $X2=0 $Y2=0
cc_289 N_A_59_463#_c_227_n N_A_688_126#_c_1080_n 0.0182498f $X=3.525 $Y=1.185
+ $X2=0 $Y2=0
cc_290 N_A_59_463#_c_232_n N_A_688_126#_c_1080_n 4.97159e-19 $X=3.795 $Y=1.715
+ $X2=0 $Y2=0
cc_291 N_A_59_463#_M1004_g N_A_688_126#_c_1083_n 0.00398235f $X=3.52 $Y=2.525
+ $X2=0 $Y2=0
cc_292 N_A_59_463#_c_229_n N_A_688_126#_c_1083_n 0.00336233f $X=3.61 $Y=1.715
+ $X2=0 $Y2=0
cc_293 N_A_59_463#_c_232_n N_A_688_126#_c_1083_n 0.00502552f $X=3.795 $Y=1.715
+ $X2=0 $Y2=0
cc_294 N_A_59_463#_M1016_g N_A_688_126#_c_1071_n 0.00716405f $X=3.795 $Y=0.84
+ $X2=0 $Y2=0
cc_295 N_A_59_463#_c_227_n N_A_688_126#_c_1071_n 0.0137765f $X=3.525 $Y=1.185
+ $X2=0 $Y2=0
cc_296 N_A_59_463#_c_229_n N_A_688_126#_c_1071_n 0.0321509f $X=3.61 $Y=1.715
+ $X2=0 $Y2=0
cc_297 N_A_59_463#_M1004_g N_A_688_126#_c_1074_n 0.00604731f $X=3.52 $Y=2.525
+ $X2=0 $Y2=0
cc_298 N_A_59_463#_c_229_n N_A_688_126#_c_1078_n 0.0119782f $X=3.61 $Y=1.715
+ $X2=0 $Y2=0
cc_299 N_A_59_463#_c_232_n N_A_688_126#_c_1078_n 0.00185768f $X=3.795 $Y=1.715
+ $X2=0 $Y2=0
cc_300 N_A_59_463#_c_220_n N_VGND_c_1145_n 0.0185118f $X=1.52 $Y=1.22 $X2=0
+ $Y2=0
cc_301 N_A_59_463#_c_221_n N_VGND_c_1145_n 0.00957848f $X=1.605 $Y=1.135 $X2=0
+ $Y2=0
cc_302 N_A_59_463#_c_225_n N_VGND_c_1145_n 0.00989869f $X=1.69 $Y=0.36 $X2=0
+ $Y2=0
cc_303 N_A_59_463#_c_224_n N_VGND_c_1146_n 0.0138929f $X=2.355 $Y=0.36 $X2=0
+ $Y2=0
cc_304 N_A_59_463#_c_226_n N_VGND_c_1146_n 0.0326123f $X=2.44 $Y=1.1 $X2=0 $Y2=0
cc_305 N_A_59_463#_c_227_n N_VGND_c_1146_n 0.0140071f $X=3.525 $Y=1.185 $X2=0
+ $Y2=0
cc_306 N_A_59_463#_c_224_n N_VGND_c_1149_n 0.0484125f $X=2.355 $Y=0.36 $X2=0
+ $Y2=0
cc_307 N_A_59_463#_c_225_n N_VGND_c_1149_n 0.0108121f $X=1.69 $Y=0.36 $X2=0
+ $Y2=0
cc_308 N_A_59_463#_M1016_g N_VGND_c_1156_n 9.43998e-19 $X=3.795 $Y=0.84 $X2=0
+ $Y2=0
cc_309 N_A_59_463#_c_224_n N_VGND_c_1156_n 0.027755f $X=2.355 $Y=0.36 $X2=0
+ $Y2=0
cc_310 N_A_59_463#_c_225_n N_VGND_c_1156_n 0.00586676f $X=1.69 $Y=0.36 $X2=0
+ $Y2=0
cc_311 N_A_59_463#_c_230_n N_VGND_c_1156_n 0.00216434f $X=0.535 $Y=0.905 $X2=0
+ $Y2=0
cc_312 N_A_59_463#_c_226_n A_453_126# 0.00349834f $X=2.44 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_313 N_A3_M1003_g N_A1_M1022_g 0.02272f $X=2.55 $Y=0.84 $X2=0 $Y2=0
cc_314 N_A3_M1007_g N_A1_M1011_g 0.0110116f $X=2.44 $Y=2.525 $X2=0 $Y2=0
cc_315 N_A3_c_361_n N_A1_c_406_n 0.0145709f $X=2.53 $Y=1.895 $X2=0 $Y2=0
cc_316 N_A3_c_366_n N_A1_c_410_n 0.0145709f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_317 A3 N_A1_c_407_n 0.00289676f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_318 N_A3_c_363_n N_A1_c_407_n 0.0145709f $X=2.53 $Y=1.555 $X2=0 $Y2=0
cc_319 A3 N_A1_c_420_n 0.0388899f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A3_c_363_n N_A1_c_420_n 5.96644e-19 $X=2.53 $Y=1.555 $X2=0 $Y2=0
cc_321 N_A3_M1007_g N_S0_c_463_n 0.0103334f $X=2.44 $Y=2.525 $X2=0 $Y2=0
cc_322 N_A3_M1003_g N_S0_M1006_g 0.0396571f $X=2.55 $Y=0.84 $X2=0 $Y2=0
cc_323 N_A3_M1003_g N_S0_c_451_n 0.008526f $X=2.55 $Y=0.84 $X2=0 $Y2=0
cc_324 N_A3_M1007_g N_VPWR_c_832_n 0.00813738f $X=2.44 $Y=2.525 $X2=0 $Y2=0
cc_325 N_A3_M1007_g N_VPWR_c_830_n 8.20269e-19 $X=2.44 $Y=2.525 $X2=0 $Y2=0
cc_326 N_A3_M1003_g N_A_345_126#_c_914_n 0.0028487f $X=2.55 $Y=0.84 $X2=0 $Y2=0
cc_327 N_A3_c_366_n N_A_345_126#_c_914_n 0.00384775f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_328 A3 N_A_345_126#_c_914_n 0.035434f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_329 N_A3_c_363_n N_A_345_126#_c_914_n 0.00352076f $X=2.53 $Y=1.555 $X2=0
+ $Y2=0
cc_330 N_A3_M1007_g N_A_345_126#_c_921_n 0.0150063f $X=2.44 $Y=2.525 $X2=0 $Y2=0
cc_331 N_A3_c_366_n N_A_345_126#_c_921_n 0.00508874f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_332 A3 N_A_345_126#_c_921_n 0.0247988f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_333 N_A3_M1007_g N_A_345_126#_c_951_n 0.00275012f $X=2.44 $Y=2.525 $X2=0
+ $Y2=0
cc_334 N_A3_M1007_g N_A_345_126#_c_924_n 2.95692e-19 $X=2.44 $Y=2.525 $X2=0
+ $Y2=0
cc_335 N_A3_M1003_g N_A_345_126#_c_919_n 2.87936e-19 $X=2.55 $Y=0.84 $X2=0 $Y2=0
cc_336 N_A3_M1003_g N_VGND_c_1146_n 0.00175725f $X=2.55 $Y=0.84 $X2=0 $Y2=0
cc_337 N_A3_M1003_g N_VGND_c_1156_n 6.31978e-19 $X=2.55 $Y=0.84 $X2=0 $Y2=0
cc_338 N_A1_M1011_g N_S0_c_463_n 0.00890008f $X=3.16 $Y=2.525 $X2=0 $Y2=0
cc_339 N_A1_M1022_g N_S0_c_451_n 0.00908269f $X=3.005 $Y=0.84 $X2=0 $Y2=0
cc_340 N_A1_M1022_g N_S0_M1015_g 0.0420433f $X=3.005 $Y=0.84 $X2=0 $Y2=0
cc_341 N_A1_M1011_g N_VPWR_c_832_n 0.00120922f $X=3.16 $Y=2.525 $X2=0 $Y2=0
cc_342 N_A1_M1011_g N_A_345_126#_c_921_n 0.00862852f $X=3.16 $Y=2.525 $X2=0
+ $Y2=0
cc_343 N_A1_c_410_n N_A_345_126#_c_921_n 0.00520455f $X=3.07 $Y=2.06 $X2=0 $Y2=0
cc_344 N_A1_c_420_n N_A_345_126#_c_921_n 0.0199025f $X=3.07 $Y=1.555 $X2=0 $Y2=0
cc_345 N_A1_M1011_g N_A_345_126#_c_951_n 0.0122675f $X=3.16 $Y=2.525 $X2=0 $Y2=0
cc_346 N_A1_M1011_g N_A_345_126#_c_923_n 0.00450121f $X=3.16 $Y=2.525 $X2=0
+ $Y2=0
cc_347 N_A1_M1011_g N_A_345_126#_c_924_n 0.00255095f $X=3.16 $Y=2.525 $X2=0
+ $Y2=0
cc_348 N_A1_M1022_g N_A_688_126#_c_1080_n 5.82953e-19 $X=3.005 $Y=0.84 $X2=0
+ $Y2=0
cc_349 N_A1_M1011_g N_A_688_126#_c_1083_n 5.44074e-19 $X=3.16 $Y=2.525 $X2=0
+ $Y2=0
cc_350 N_A1_c_420_n N_A_688_126#_c_1074_n 0.00229766f $X=3.07 $Y=1.555 $X2=0
+ $Y2=0
cc_351 N_A1_c_420_n N_A_688_126#_c_1078_n 4.48212e-19 $X=3.07 $Y=1.555 $X2=0
+ $Y2=0
cc_352 N_A1_M1022_g N_VGND_c_1146_n 0.00327423f $X=3.005 $Y=0.84 $X2=0 $Y2=0
cc_353 N_A1_M1022_g N_VGND_c_1156_n 9.43998e-19 $X=3.005 $Y=0.84 $X2=0 $Y2=0
cc_354 N_S0_c_453_n N_A0_c_582_n 0.00908269f $X=4.86 $Y=0.185 $X2=-0.19
+ $Y2=-0.245
cc_355 N_S0_c_454_n N_A0_c_582_n 0.00818553f $X=4.935 $Y=3.075 $X2=-0.19
+ $Y2=-0.245
cc_356 N_S0_M1017_g N_A0_M1019_g 0.0428137f $X=3.95 $Y=2.525 $X2=0 $Y2=0
cc_357 N_S0_c_466_n N_A0_M1019_g 0.00889584f $X=4.86 $Y=3.15 $X2=0 $Y2=0
cc_358 N_S0_c_454_n N_A0_M1019_g 0.031994f $X=4.935 $Y=3.075 $X2=0 $Y2=0
cc_359 N_S0_c_454_n A0 0.00339015f $X=4.935 $Y=3.075 $X2=0 $Y2=0
cc_360 N_S0_c_454_n N_A0_c_585_n 0.0126958f $X=4.935 $Y=3.075 $X2=0 $Y2=0
cc_361 N_S0_c_454_n N_A_1118_37#_c_616_n 9.55488e-19 $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_362 N_S0_c_453_n N_A_1118_37#_c_617_n 0.00688101f $X=4.86 $Y=0.185 $X2=0
+ $Y2=0
cc_363 N_S0_M1023_g N_VPWR_c_831_n 0.00359426f $X=0.635 $Y=2.525 $X2=0 $Y2=0
cc_364 N_S0_M1000_g N_VPWR_c_831_n 0.00657855f $X=1.65 $Y=2.525 $X2=0 $Y2=0
cc_365 N_S0_c_463_n N_VPWR_c_832_n 0.0255122f $X=3.875 $Y=3.15 $X2=0 $Y2=0
cc_366 N_S0_M1017_g N_VPWR_c_833_n 0.0038758f $X=3.95 $Y=2.525 $X2=0 $Y2=0
cc_367 N_S0_c_466_n N_VPWR_c_833_n 0.0165604f $X=4.86 $Y=3.15 $X2=0 $Y2=0
cc_368 N_S0_c_454_n N_VPWR_c_833_n 0.00632963f $X=4.935 $Y=3.075 $X2=0 $Y2=0
cc_369 N_S0_M1023_g N_VPWR_c_835_n 0.00431487f $X=0.635 $Y=2.525 $X2=0 $Y2=0
cc_370 N_S0_c_463_n N_VPWR_c_837_n 0.0447285f $X=3.875 $Y=3.15 $X2=0 $Y2=0
cc_371 N_S0_c_464_n N_VPWR_c_839_n 0.0308935f $X=1.725 $Y=3.15 $X2=0 $Y2=0
cc_372 N_S0_c_466_n N_VPWR_c_840_n 0.0090328f $X=4.86 $Y=3.15 $X2=0 $Y2=0
cc_373 N_S0_M1023_g N_VPWR_c_830_n 0.00477801f $X=0.635 $Y=2.525 $X2=0 $Y2=0
cc_374 N_S0_c_463_n N_VPWR_c_830_n 0.060014f $X=3.875 $Y=3.15 $X2=0 $Y2=0
cc_375 N_S0_c_464_n N_VPWR_c_830_n 0.0116041f $X=1.725 $Y=3.15 $X2=0 $Y2=0
cc_376 N_S0_c_466_n N_VPWR_c_830_n 0.033744f $X=4.86 $Y=3.15 $X2=0 $Y2=0
cc_377 N_S0_c_468_n N_VPWR_c_830_n 0.00385141f $X=3.95 $Y=3.15 $X2=0 $Y2=0
cc_378 N_S0_c_463_n N_A_345_126#_c_974_n 0.00299556f $X=3.875 $Y=3.15 $X2=0
+ $Y2=0
cc_379 N_S0_M1006_g N_A_345_126#_c_914_n 0.00583334f $X=2.19 $Y=0.84 $X2=0 $Y2=0
cc_380 N_S0_M1000_g N_A_345_126#_c_922_n 0.00183973f $X=1.65 $Y=2.525 $X2=0
+ $Y2=0
cc_381 N_S0_c_463_n N_A_345_126#_c_923_n 0.00985759f $X=3.875 $Y=3.15 $X2=0
+ $Y2=0
cc_382 N_S0_M1017_g N_A_345_126#_c_923_n 0.0114249f $X=3.95 $Y=2.525 $X2=0 $Y2=0
cc_383 N_S0_c_466_n N_A_345_126#_c_923_n 0.00402004f $X=4.86 $Y=3.15 $X2=0 $Y2=0
cc_384 N_S0_c_463_n N_A_345_126#_c_924_n 0.00256652f $X=3.875 $Y=3.15 $X2=0
+ $Y2=0
cc_385 N_S0_M1017_g N_A_345_126#_c_925_n 9.34571e-19 $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_386 N_S0_c_454_n N_A_345_126#_c_925_n 8.11741e-19 $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_387 N_S0_c_454_n N_A_345_126#_c_926_n 0.0129418f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_388 N_S0_M1017_g N_A_345_126#_c_927_n 2.21919e-19 $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_389 N_S0_c_454_n N_A_345_126#_c_928_n 0.0184326f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_390 N_S0_c_454_n N_A_345_126#_c_930_n 0.00773309f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_391 N_S0_c_454_n N_A_345_126#_c_915_n 0.00679002f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_392 N_S0_c_454_n N_A_345_126#_c_917_n 0.00440591f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_393 N_S0_M1006_g N_A_345_126#_c_919_n 0.00518141f $X=2.19 $Y=0.84 $X2=0 $Y2=0
cc_394 N_S0_M1015_g N_A_688_126#_c_1080_n 0.00446994f $X=3.365 $Y=0.84 $X2=0
+ $Y2=0
cc_395 N_S0_c_453_n N_A_688_126#_c_1080_n 0.00604501f $X=4.86 $Y=0.185 $X2=0
+ $Y2=0
cc_396 N_S0_M1017_g N_A_688_126#_c_1083_n 0.00553673f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_397 N_S0_M1017_g N_A_688_126#_c_1074_n 0.00807192f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_398 N_S0_c_454_n N_A_688_126#_c_1075_n 0.0176611f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_399 N_S0_c_454_n N_A_688_126#_c_1072_n 0.0208658f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_400 N_S0_c_454_n N_A_688_126#_c_1077_n 0.00868914f $X=4.935 $Y=3.075 $X2=0
+ $Y2=0
cc_401 N_S0_c_449_n N_VGND_c_1145_n 0.0252521f $X=2.115 $Y=0.185 $X2=0 $Y2=0
cc_402 N_S0_c_458_n N_VGND_c_1145_n 0.0116505f $X=0.51 $Y=0.35 $X2=0 $Y2=0
cc_403 N_S0_c_459_n N_VGND_c_1145_n 0.0106453f $X=0.585 $Y=0.185 $X2=0 $Y2=0
cc_404 N_S0_c_460_n N_VGND_c_1145_n 0.00694768f $X=0.24 $Y=0.35 $X2=0 $Y2=0
cc_405 N_S0_M1006_g N_VGND_c_1146_n 0.0011604f $X=2.19 $Y=0.84 $X2=0 $Y2=0
cc_406 N_S0_c_451_n N_VGND_c_1146_n 0.0183639f $X=3.29 $Y=0.185 $X2=0 $Y2=0
cc_407 N_S0_M1015_g N_VGND_c_1146_n 0.00725446f $X=3.365 $Y=0.84 $X2=0 $Y2=0
cc_408 N_S0_c_453_n N_VGND_c_1147_n 0.0193554f $X=4.86 $Y=0.185 $X2=0 $Y2=0
cc_409 N_S0_c_454_n N_VGND_c_1147_n 0.0125586f $X=4.935 $Y=3.075 $X2=0 $Y2=0
cc_410 N_S0_c_449_n N_VGND_c_1149_n 0.0385976f $X=2.115 $Y=0.185 $X2=0 $Y2=0
cc_411 N_S0_c_451_n N_VGND_c_1151_n 0.0428273f $X=3.29 $Y=0.185 $X2=0 $Y2=0
cc_412 N_S0_c_458_n N_VGND_c_1153_n 0.0202769f $X=0.51 $Y=0.35 $X2=0 $Y2=0
cc_413 N_S0_c_459_n N_VGND_c_1153_n 0.0152618f $X=0.585 $Y=0.185 $X2=0 $Y2=0
cc_414 N_S0_c_460_n N_VGND_c_1153_n 0.0108395f $X=0.24 $Y=0.35 $X2=0 $Y2=0
cc_415 N_S0_c_453_n N_VGND_c_1154_n 0.0195671f $X=4.86 $Y=0.185 $X2=0 $Y2=0
cc_416 N_S0_c_449_n N_VGND_c_1156_n 0.0306959f $X=2.115 $Y=0.185 $X2=0 $Y2=0
cc_417 N_S0_c_451_n N_VGND_c_1156_n 0.032289f $X=3.29 $Y=0.185 $X2=0 $Y2=0
cc_418 N_S0_c_453_n N_VGND_c_1156_n 0.0580698f $X=4.86 $Y=0.185 $X2=0 $Y2=0
cc_419 N_S0_c_456_n N_VGND_c_1156_n 0.00371918f $X=2.19 $Y=0.185 $X2=0 $Y2=0
cc_420 N_S0_c_457_n N_VGND_c_1156_n 0.00847832f $X=3.365 $Y=0.185 $X2=0 $Y2=0
cc_421 N_S0_c_458_n N_VGND_c_1156_n 0.0115698f $X=0.51 $Y=0.35 $X2=0 $Y2=0
cc_422 N_S0_c_459_n N_VGND_c_1156_n 0.0179593f $X=0.585 $Y=0.185 $X2=0 $Y2=0
cc_423 N_S0_c_460_n N_VGND_c_1156_n 0.00640038f $X=0.24 $Y=0.35 $X2=0 $Y2=0
cc_424 N_A0_M1019_g N_VPWR_c_833_n 0.00160775f $X=4.31 $Y=2.525 $X2=0 $Y2=0
cc_425 N_A0_M1019_g N_A_345_126#_c_923_n 0.00402945f $X=4.31 $Y=2.525 $X2=0
+ $Y2=0
cc_426 N_A0_M1019_g N_A_345_126#_c_925_n 0.0111803f $X=4.31 $Y=2.525 $X2=0 $Y2=0
cc_427 N_A0_M1019_g N_A_345_126#_c_927_n 0.00864472f $X=4.31 $Y=2.525 $X2=0
+ $Y2=0
cc_428 N_A0_M1019_g N_A_345_126#_c_928_n 2.80284e-19 $X=4.31 $Y=2.525 $X2=0
+ $Y2=0
cc_429 N_A0_c_582_n N_A_688_126#_c_1071_n 0.00433825f $X=4.155 $Y=1.16 $X2=0
+ $Y2=0
cc_430 A0 N_A_688_126#_c_1071_n 0.0174988f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_431 N_A0_c_585_n N_A_688_126#_c_1071_n 0.00638479f $X=4.31 $Y=1.325 $X2=0
+ $Y2=0
cc_432 N_A0_M1019_g N_A_688_126#_c_1074_n 0.0050458f $X=4.31 $Y=2.525 $X2=0
+ $Y2=0
cc_433 N_A0_M1019_g N_A_688_126#_c_1075_n 0.0141243f $X=4.31 $Y=2.525 $X2=0
+ $Y2=0
cc_434 A0 N_A_688_126#_c_1075_n 0.0195361f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_435 N_A0_c_585_n N_A_688_126#_c_1075_n 0.00880049f $X=4.31 $Y=1.325 $X2=0
+ $Y2=0
cc_436 A0 N_A_688_126#_c_1072_n 0.0105188f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_437 N_A0_c_582_n N_VGND_c_1147_n 0.0038288f $X=4.155 $Y=1.16 $X2=0 $Y2=0
cc_438 A0 N_VGND_c_1147_n 0.0107638f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_439 N_A0_c_585_n N_VGND_c_1147_n 0.00563489f $X=4.31 $Y=1.325 $X2=0 $Y2=0
cc_440 N_A0_c_582_n N_VGND_c_1156_n 9.43998e-19 $X=4.155 $Y=1.16 $X2=0 $Y2=0
cc_441 N_A_1118_37#_c_619_n N_S1_M1012_g 0.0106605f $X=5.92 $Y=1.87 $X2=0 $Y2=0
cc_442 N_A_1118_37#_M1005_g N_S1_M1012_g 0.0133934f $X=6.275 $Y=2.525 $X2=0
+ $Y2=0
cc_443 N_A_1118_37#_M1005_g N_S1_c_694_n 0.00883541f $X=6.275 $Y=2.525 $X2=0
+ $Y2=0
cc_444 N_A_1118_37#_M1018_g N_S1_c_685_n 0.0186138f $X=5.845 $Y=1.065 $X2=0
+ $Y2=0
cc_445 N_A_1118_37#_c_616_n N_S1_c_685_n 7.86069e-19 $X=6.935 $Y=0.35 $X2=0
+ $Y2=0
cc_446 N_A_1118_37#_c_622_n N_S1_c_687_n 0.0213055f $X=6.51 $Y=1.97 $X2=0 $Y2=0
cc_447 N_A_1118_37#_c_623_n N_S1_c_696_n 0.00401349f $X=7.04 $Y=2.78 $X2=0 $Y2=0
cc_448 N_A_1118_37#_M1005_g N_S1_c_688_n 0.00198571f $X=6.275 $Y=2.525 $X2=0
+ $Y2=0
cc_449 N_A_1118_37#_c_621_n N_S1_c_688_n 0.00799933f $X=6.935 $Y=1.97 $X2=0
+ $Y2=0
cc_450 N_A_1118_37#_c_622_n N_S1_c_688_n 0.0152222f $X=6.51 $Y=1.97 $X2=0 $Y2=0
cc_451 N_A_1118_37#_c_623_n N_S1_c_688_n 0.00807867f $X=7.04 $Y=2.78 $X2=0 $Y2=0
cc_452 N_A_1118_37#_c_623_n N_S1_c_698_n 0.00159169f $X=7.04 $Y=2.78 $X2=0 $Y2=0
cc_453 N_A_1118_37#_M1005_g N_S1_c_699_n 0.00948828f $X=6.275 $Y=2.525 $X2=0
+ $Y2=0
cc_454 N_A_1118_37#_c_621_n N_S1_c_699_n 0.00861993f $X=6.935 $Y=1.97 $X2=0
+ $Y2=0
cc_455 N_A_1118_37#_c_623_n N_S1_c_699_n 0.0127725f $X=7.04 $Y=2.78 $X2=0 $Y2=0
cc_456 N_A_1118_37#_c_616_n N_S1_c_690_n 0.00335802f $X=6.935 $Y=0.35 $X2=0
+ $Y2=0
cc_457 N_A_1118_37#_c_643_p N_S1_c_690_n 0.00555802f $X=7.04 $Y=0.35 $X2=0 $Y2=0
cc_458 N_A_1118_37#_c_616_n S1 0.00484322f $X=6.935 $Y=0.35 $X2=0 $Y2=0
cc_459 N_A_1118_37#_c_643_p S1 0.0107536f $X=7.04 $Y=0.35 $X2=0 $Y2=0
cc_460 N_A_1118_37#_c_621_n N_A_1184_171#_M1002_g 0.00153007f $X=6.935 $Y=1.97
+ $X2=0 $Y2=0
cc_461 N_A_1118_37#_c_623_n N_A_1184_171#_M1002_g 0.00365613f $X=7.04 $Y=2.78
+ $X2=0 $Y2=0
cc_462 N_A_1118_37#_M1018_g N_A_1184_171#_c_771_n 0.00186917f $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_463 N_A_1118_37#_M1018_g N_A_1184_171#_c_778_n 0.00197212f $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_464 N_A_1118_37#_c_621_n N_A_1184_171#_c_778_n 0.0127311f $X=6.935 $Y=1.97
+ $X2=0 $Y2=0
cc_465 N_A_1118_37#_c_622_n N_A_1184_171#_c_778_n 0.0120698f $X=6.51 $Y=1.97
+ $X2=0 $Y2=0
cc_466 N_A_1118_37#_c_624_n N_A_1184_171#_c_778_n 0.0184546f $X=6.2 $Y=1.965
+ $X2=0 $Y2=0
cc_467 N_A_1118_37#_c_621_n N_A_1184_171#_c_772_n 0.0571537f $X=6.935 $Y=1.97
+ $X2=0 $Y2=0
cc_468 N_A_1118_37#_c_624_n N_A_1184_171#_c_772_n 0.00713363f $X=6.2 $Y=1.965
+ $X2=0 $Y2=0
cc_469 N_A_1118_37#_M1018_g N_A_1184_171#_c_775_n 0.00395151f $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_470 N_A_1118_37#_c_623_n N_VPWR_c_840_n 0.0075246f $X=7.04 $Y=2.78 $X2=0
+ $Y2=0
cc_471 N_A_1118_37#_c_623_n N_VPWR_c_830_n 0.00751788f $X=7.04 $Y=2.78 $X2=0
+ $Y2=0
cc_472 N_A_1118_37#_M1018_g N_A_345_126#_c_915_n 0.0294719f $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_473 N_A_1118_37#_c_619_n N_A_345_126#_c_915_n 0.00528896f $X=5.92 $Y=1.87
+ $X2=0 $Y2=0
cc_474 N_A_1118_37#_M1005_g N_A_345_126#_c_915_n 6.13421e-19 $X=6.275 $Y=2.525
+ $X2=0 $Y2=0
cc_475 N_A_1118_37#_M1018_g N_A_345_126#_c_916_n 0.0124391f $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_476 N_A_1118_37#_c_616_n N_A_345_126#_c_916_n 0.0546684f $X=6.935 $Y=0.35
+ $X2=0 $Y2=0
cc_477 N_A_1118_37#_M1018_g N_A_345_126#_c_917_n 0.00370163f $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_478 N_A_1118_37#_c_616_n N_A_345_126#_c_917_n 0.0120962f $X=6.935 $Y=0.35
+ $X2=0 $Y2=0
cc_479 N_A_1118_37#_c_617_n N_A_345_126#_c_917_n 0.00370505f $X=5.755 $Y=0.35
+ $X2=0 $Y2=0
cc_480 N_A_1118_37#_M1005_g N_A_345_126#_c_932_n 0.00948176f $X=6.275 $Y=2.525
+ $X2=0 $Y2=0
cc_481 N_A_1118_37#_c_622_n N_A_345_126#_c_932_n 7.7796e-19 $X=6.51 $Y=1.97
+ $X2=0 $Y2=0
cc_482 N_A_1118_37#_c_623_n N_A_345_126#_c_932_n 0.00717777f $X=7.04 $Y=2.78
+ $X2=0 $Y2=0
cc_483 N_A_1118_37#_M1005_g N_A_345_126#_c_933_n 9.58968e-19 $X=6.275 $Y=2.525
+ $X2=0 $Y2=0
cc_484 N_A_1118_37#_c_621_n N_A_345_126#_c_933_n 0.0083602f $X=6.935 $Y=1.97
+ $X2=0 $Y2=0
cc_485 N_A_1118_37#_c_622_n N_A_345_126#_c_933_n 0.00459042f $X=6.51 $Y=1.97
+ $X2=0 $Y2=0
cc_486 N_A_1118_37#_c_623_n N_A_345_126#_c_933_n 0.0171021f $X=7.04 $Y=2.78
+ $X2=0 $Y2=0
cc_487 N_A_1118_37#_M1018_g N_A_688_126#_c_1072_n 0.00382288f $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_488 N_A_1118_37#_c_619_n N_A_688_126#_c_1077_n 2.41375e-19 $X=5.92 $Y=1.87
+ $X2=0 $Y2=0
cc_489 N_A_1118_37#_M1018_g N_A_688_126#_c_1079_n 9.46911e-19 $X=5.845 $Y=1.065
+ $X2=0 $Y2=0
cc_490 N_A_1118_37#_c_621_n N_X_c_1132_n 0.00563618f $X=6.935 $Y=1.97 $X2=0
+ $Y2=0
cc_491 N_A_1118_37#_c_623_n N_X_c_1132_n 0.0168489f $X=7.04 $Y=2.78 $X2=0 $Y2=0
cc_492 N_A_1118_37#_c_616_n N_VGND_c_1154_n 0.0805878f $X=6.935 $Y=0.35 $X2=0
+ $Y2=0
cc_493 N_A_1118_37#_c_617_n N_VGND_c_1154_n 0.00651318f $X=5.755 $Y=0.35 $X2=0
+ $Y2=0
cc_494 N_A_1118_37#_c_643_p N_VGND_c_1154_n 0.0124385f $X=7.04 $Y=0.35 $X2=0
+ $Y2=0
cc_495 N_A_1118_37#_M1025_s N_VGND_c_1156_n 0.00255657f $X=6.915 $Y=0.235 $X2=0
+ $Y2=0
cc_496 N_A_1118_37#_c_616_n N_VGND_c_1156_n 0.0487561f $X=6.935 $Y=0.35 $X2=0
+ $Y2=0
cc_497 N_A_1118_37#_c_617_n N_VGND_c_1156_n 0.00976432f $X=5.755 $Y=0.35 $X2=0
+ $Y2=0
cc_498 N_A_1118_37#_c_643_p N_VGND_c_1156_n 0.00789949f $X=7.04 $Y=0.35 $X2=0
+ $Y2=0
cc_499 N_S1_c_691_n N_A_1184_171#_c_769_n 0.0127994f $X=6.96 $Y=1.46 $X2=0 $Y2=0
cc_500 N_S1_c_689_n N_A_1184_171#_M1008_g 0.0224564f $X=7.255 $Y=0.765 $X2=0
+ $Y2=0
cc_501 S1 N_A_1184_171#_M1008_g 0.00207005f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_502 N_S1_c_692_n N_A_1184_171#_M1008_g 0.00407663f $X=6.96 $Y=0.93 $X2=0
+ $Y2=0
cc_503 N_S1_c_688_n N_A_1184_171#_M1002_g 0.00855433f $X=7.05 $Y=2.375 $X2=0
+ $Y2=0
cc_504 N_S1_c_699_n N_A_1184_171#_M1002_g 0.0209497f $X=7.255 $Y=2.45 $X2=0
+ $Y2=0
cc_505 N_S1_c_685_n N_A_1184_171#_c_771_n 0.00582002f $X=6.275 $Y=1.385 $X2=0
+ $Y2=0
cc_506 S1 N_A_1184_171#_c_771_n 0.00359104f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_507 N_S1_M1012_g N_A_1184_171#_c_778_n 9.34584e-19 $X=5.845 $Y=2.525 $X2=0
+ $Y2=0
cc_508 N_S1_c_687_n N_A_1184_171#_c_772_n 0.0209698f $X=6.35 $Y=1.46 $X2=0 $Y2=0
cc_509 N_S1_c_688_n N_A_1184_171#_c_772_n 0.0102115f $X=7.05 $Y=2.375 $X2=0
+ $Y2=0
cc_510 N_S1_c_699_n N_A_1184_171#_c_772_n 0.00500174f $X=7.255 $Y=2.45 $X2=0
+ $Y2=0
cc_511 N_S1_c_690_n N_A_1184_171#_c_772_n 0.00508767f $X=7.255 $Y=0.84 $X2=0
+ $Y2=0
cc_512 S1 N_A_1184_171#_c_772_n 0.023986f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_513 N_S1_c_688_n N_A_1184_171#_c_780_n 8.51393e-19 $X=7.05 $Y=2.375 $X2=0
+ $Y2=0
cc_514 S1 N_A_1184_171#_c_773_n 0.00710126f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_515 N_S1_c_692_n N_A_1184_171#_c_773_n 0.00167108f $X=6.96 $Y=0.93 $X2=0
+ $Y2=0
cc_516 S1 N_A_1184_171#_c_774_n 6.59556e-19 $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_517 N_S1_c_692_n N_A_1184_171#_c_774_n 0.0127994f $X=6.96 $Y=0.93 $X2=0 $Y2=0
cc_518 N_S1_c_688_n N_A_1184_171#_c_782_n 0.0127994f $X=7.05 $Y=2.375 $X2=0
+ $Y2=0
cc_519 N_S1_c_696_n N_VPWR_c_834_n 0.0011069f $X=6.765 $Y=3.075 $X2=0 $Y2=0
cc_520 N_S1_c_698_n N_VPWR_c_834_n 0.00290284f $X=7.255 $Y=2.525 $X2=0 $Y2=0
cc_521 N_S1_c_695_n N_VPWR_c_840_n 0.0281018f $X=5.92 $Y=3.15 $X2=0 $Y2=0
cc_522 N_S1_c_698_n N_VPWR_c_840_n 0.00545548f $X=7.255 $Y=2.525 $X2=0 $Y2=0
cc_523 N_S1_c_694_n N_VPWR_c_830_n 0.0325052f $X=6.69 $Y=3.15 $X2=0 $Y2=0
cc_524 N_S1_c_695_n N_VPWR_c_830_n 0.0061073f $X=5.92 $Y=3.15 $X2=0 $Y2=0
cc_525 N_S1_c_698_n N_VPWR_c_830_n 0.0104976f $X=7.255 $Y=2.525 $X2=0 $Y2=0
cc_526 N_S1_M1012_g N_A_345_126#_c_928_n 0.00113093f $X=5.845 $Y=2.525 $X2=0
+ $Y2=0
cc_527 N_S1_M1012_g N_A_345_126#_c_915_n 0.0188167f $X=5.845 $Y=2.525 $X2=0
+ $Y2=0
cc_528 N_S1_c_685_n N_A_345_126#_c_915_n 6.52871e-19 $X=6.275 $Y=1.385 $X2=0
+ $Y2=0
cc_529 N_S1_c_685_n N_A_345_126#_c_916_n 0.0116343f $X=6.275 $Y=1.385 $X2=0
+ $Y2=0
cc_530 N_S1_c_689_n N_A_345_126#_c_916_n 0.00388418f $X=7.255 $Y=0.765 $X2=0
+ $Y2=0
cc_531 N_S1_c_690_n N_A_345_126#_c_916_n 5.94742e-19 $X=7.255 $Y=0.84 $X2=0
+ $Y2=0
cc_532 N_S1_M1012_g N_A_345_126#_c_932_n 0.0121191f $X=5.845 $Y=2.525 $X2=0
+ $Y2=0
cc_533 N_S1_c_694_n N_A_345_126#_c_932_n 0.0108713f $X=6.69 $Y=3.15 $X2=0 $Y2=0
cc_534 N_S1_c_696_n N_A_345_126#_c_932_n 0.00400676f $X=6.765 $Y=3.075 $X2=0
+ $Y2=0
cc_535 N_S1_c_685_n N_A_345_126#_c_918_n 0.00105038f $X=6.275 $Y=1.385 $X2=0
+ $Y2=0
cc_536 N_S1_c_686_n N_A_345_126#_c_918_n 0.00327544f $X=6.795 $Y=1.46 $X2=0
+ $Y2=0
cc_537 N_S1_c_690_n N_A_345_126#_c_918_n 0.00409379f $X=7.255 $Y=0.84 $X2=0
+ $Y2=0
cc_538 S1 N_A_345_126#_c_918_n 0.0214957f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_539 N_S1_c_699_n N_A_345_126#_c_933_n 0.00380769f $X=7.255 $Y=2.45 $X2=0
+ $Y2=0
cc_540 N_S1_M1012_g N_A_345_126#_c_934_n 0.00480547f $X=5.845 $Y=2.525 $X2=0
+ $Y2=0
cc_541 N_S1_M1012_g N_A_688_126#_c_1077_n 0.00219462f $X=5.845 $Y=2.525 $X2=0
+ $Y2=0
cc_542 S1 N_X_c_1132_n 0.0092641f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_543 N_S1_c_689_n N_VGND_c_1148_n 0.00274937f $X=7.255 $Y=0.765 $X2=0 $Y2=0
cc_544 N_S1_c_689_n N_VGND_c_1154_n 0.00585385f $X=7.255 $Y=0.765 $X2=0 $Y2=0
cc_545 N_S1_c_690_n N_VGND_c_1154_n 7.55273e-19 $X=7.255 $Y=0.84 $X2=0 $Y2=0
cc_546 N_S1_c_689_n N_VGND_c_1156_n 0.0119704f $X=7.255 $Y=0.765 $X2=0 $Y2=0
cc_547 N_S1_c_690_n N_VGND_c_1156_n 7.80545e-19 $X=7.255 $Y=0.84 $X2=0 $Y2=0
cc_548 S1 N_VGND_c_1156_n 8.39253e-19 $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_549 N_A_1184_171#_M1002_g N_VPWR_c_834_n 0.00290284f $X=7.685 $Y=2.845 $X2=0
+ $Y2=0
cc_550 N_A_1184_171#_M1002_g N_VPWR_c_841_n 0.00545548f $X=7.685 $Y=2.845 $X2=0
+ $Y2=0
cc_551 N_A_1184_171#_M1002_g N_VPWR_c_830_n 0.0111011f $X=7.685 $Y=2.845 $X2=0
+ $Y2=0
cc_552 N_A_1184_171#_c_771_n N_A_345_126#_c_915_n 0.0279338f $X=6.06 $Y=1.13
+ $X2=0 $Y2=0
cc_553 N_A_1184_171#_c_778_n N_A_345_126#_c_915_n 0.0524381f $X=6.06 $Y=2.46
+ $X2=0 $Y2=0
cc_554 N_A_1184_171#_c_775_n N_A_345_126#_c_915_n 0.0131377f $X=6.07 $Y=1.62
+ $X2=0 $Y2=0
cc_555 N_A_1184_171#_c_771_n N_A_345_126#_c_916_n 0.0139641f $X=6.06 $Y=1.13
+ $X2=0 $Y2=0
cc_556 N_A_1184_171#_c_778_n N_A_345_126#_c_932_n 0.0133017f $X=6.06 $Y=2.46
+ $X2=0 $Y2=0
cc_557 N_A_1184_171#_c_772_n N_A_345_126#_c_918_n 0.00913841f $X=7.445 $Y=1.62
+ $X2=0 $Y2=0
cc_558 N_A_1184_171#_M1008_g N_X_c_1132_n 0.0588948f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_559 N_A_1184_171#_c_780_n N_X_c_1132_n 0.0240219f $X=7.53 $Y=1.535 $X2=0
+ $Y2=0
cc_560 N_A_1184_171#_c_773_n N_X_c_1132_n 0.0239766f $X=7.53 $Y=1.355 $X2=0
+ $Y2=0
cc_561 N_A_1184_171#_M1008_g N_VGND_c_1148_n 0.00285763f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_562 N_A_1184_171#_c_773_n N_VGND_c_1148_n 0.00350934f $X=7.53 $Y=1.355 $X2=0
+ $Y2=0
cc_563 N_A_1184_171#_c_774_n N_VGND_c_1148_n 0.00239796f $X=7.53 $Y=1.355 $X2=0
+ $Y2=0
cc_564 N_A_1184_171#_M1008_g N_VGND_c_1155_n 0.00585385f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_565 N_A_1184_171#_M1008_g N_VGND_c_1156_n 0.0117282f $X=7.685 $Y=0.445 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_832_n N_A_345_126#_c_974_n 0.00347818f $X=2.66 $Y=2.61 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_839_n N_A_345_126#_c_974_n 0.00322187f $X=2.495 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_830_n N_A_345_126#_c_974_n 0.00577667f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_569 N_VPWR_M1007_d N_A_345_126#_c_921_n 0.00994894f $X=2.515 $Y=2.315 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_832_n N_A_345_126#_c_921_n 0.0209862f $X=2.66 $Y=2.61 $X2=0
+ $Y2=0
cc_571 N_VPWR_M1007_d N_A_345_126#_c_951_n 0.0047605f $X=2.515 $Y=2.315 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_832_n N_A_345_126#_c_951_n 0.016106f $X=2.66 $Y=2.61 $X2=0 $Y2=0
cc_573 N_VPWR_c_833_n N_A_345_126#_c_923_n 0.0137858f $X=4.66 $Y=2.59 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_837_n N_A_345_126#_c_923_n 0.039217f $X=4.575 $Y=3.33 $X2=0
+ $Y2=0
cc_575 N_VPWR_c_830_n N_A_345_126#_c_923_n 0.0363984f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_832_n N_A_345_126#_c_924_n 0.0144397f $X=2.66 $Y=2.61 $X2=0
+ $Y2=0
cc_577 N_VPWR_c_837_n N_A_345_126#_c_924_n 0.0060012f $X=4.575 $Y=3.33 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_830_n N_A_345_126#_c_924_n 0.00534497f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_833_n N_A_345_126#_c_925_n 0.0114401f $X=4.66 $Y=2.59 $X2=0
+ $Y2=0
cc_580 N_VPWR_c_833_n N_A_345_126#_c_926_n 0.013324f $X=4.66 $Y=2.59 $X2=0 $Y2=0
cc_581 N_VPWR_c_833_n N_A_345_126#_c_928_n 0.0255877f $X=4.66 $Y=2.59 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_840_n N_A_345_126#_c_929_n 0.0209327f $X=7.365 $Y=3.33 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_830_n N_A_345_126#_c_929_n 0.018667f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_584 N_VPWR_c_833_n N_A_345_126#_c_930_n 0.0130064f $X=4.66 $Y=2.59 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_840_n N_A_345_126#_c_930_n 0.00718429f $X=7.365 $Y=3.33 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_830_n N_A_345_126#_c_930_n 0.00584888f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_840_n N_A_345_126#_c_932_n 0.0320314f $X=7.365 $Y=3.33 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_830_n N_A_345_126#_c_932_n 0.0251295f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_840_n N_A_345_126#_c_934_n 0.00732267f $X=7.365 $Y=3.33 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_830_n N_A_345_126#_c_934_n 0.00612665f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_591 N_VPWR_c_841_n N_X_c_1132_n 0.0075246f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_592 N_VPWR_c_830_n N_X_c_1132_n 0.00751788f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_593 N_A_345_126#_c_921_n A_431_463# 0.00366293f $X=3.005 $Y=2.26 $X2=-0.19
+ $Y2=-0.245
cc_594 N_A_345_126#_c_915_n N_A_688_126#_M1018_s 0.00496803f $X=5.71 $Y=2.805
+ $X2=0 $Y2=0
cc_595 N_A_345_126#_c_915_n N_A_688_126#_M1012_s 0.00476592f $X=5.71 $Y=2.805
+ $X2=0 $Y2=0
cc_596 N_A_345_126#_c_951_n N_A_688_126#_c_1083_n 0.00777759f $X=3.09 $Y=2.745
+ $X2=0 $Y2=0
cc_597 N_A_345_126#_c_923_n N_A_688_126#_c_1083_n 0.028296f $X=4.225 $Y=2.83
+ $X2=0 $Y2=0
cc_598 N_A_345_126#_c_925_n N_A_688_126#_c_1074_n 0.00495237f $X=4.31 $Y=2.745
+ $X2=0 $Y2=0
cc_599 N_A_345_126#_c_927_n N_A_688_126#_c_1074_n 0.0137841f $X=4.395 $Y=2.16
+ $X2=0 $Y2=0
cc_600 N_A_345_126#_c_926_n N_A_688_126#_c_1075_n 0.0508492f $X=4.925 $Y=2.16
+ $X2=0 $Y2=0
cc_601 N_A_345_126#_c_927_n N_A_688_126#_c_1075_n 0.0125335f $X=4.395 $Y=2.16
+ $X2=0 $Y2=0
cc_602 N_A_345_126#_c_915_n N_A_688_126#_c_1072_n 0.0545469f $X=5.71 $Y=2.805
+ $X2=0 $Y2=0
cc_603 N_A_345_126#_c_926_n N_A_688_126#_c_1077_n 0.0137864f $X=4.925 $Y=2.16
+ $X2=0 $Y2=0
cc_604 N_A_345_126#_c_928_n N_A_688_126#_c_1077_n 0.0270265f $X=5.01 $Y=2.805
+ $X2=0 $Y2=0
cc_605 N_A_345_126#_c_929_n N_A_688_126#_c_1077_n 0.0126536f $X=5.625 $Y=2.89
+ $X2=0 $Y2=0
cc_606 N_A_345_126#_c_915_n N_A_688_126#_c_1077_n 0.05192f $X=5.71 $Y=2.805
+ $X2=0 $Y2=0
cc_607 N_A_345_126#_c_915_n N_A_688_126#_c_1079_n 0.0137868f $X=5.71 $Y=2.805
+ $X2=0 $Y2=0
cc_608 N_A_688_126#_c_1080_n N_VGND_c_1151_n 0.00808338f $X=3.875 $Y=0.815 $X2=0
+ $Y2=0
cc_609 N_A_688_126#_c_1080_n N_VGND_c_1156_n 0.0146974f $X=3.875 $Y=0.815 $X2=0
+ $Y2=0
cc_610 N_A_688_126#_c_1080_n A_774_126# 0.00153824f $X=3.875 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_611 N_X_c_1132_n N_VGND_c_1155_n 0.00877924f $X=7.9 $Y=0.51 $X2=0 $Y2=0
cc_612 N_X_M1008_d N_VGND_c_1156_n 0.0042053f $X=7.76 $Y=0.235 $X2=0 $Y2=0
cc_613 N_X_c_1132_n N_VGND_c_1156_n 0.00770513f $X=7.9 $Y=0.51 $X2=0 $Y2=0
