* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4_m A B C D VGND VNB VPB VPWR X
X0 a_116_397# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_343_397# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_116_397# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_116_397# D a_199_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND D a_116_397# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_199_397# C a_271_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_271_397# B a_343_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_116_397# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_116_397# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND B a_116_397# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
