* NGSPICE file created from sky130_fd_sc_lp__a22o_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a22o_lp A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_137_409# B1 a_243_409# VPB phighvt w=1e+06u l=250000u
+  ad=5.6e+11p pd=5.12e+06u as=5.85e+11p ps=3.17e+06u
M1001 VGND A2 a_389_47# VNB nshort w=420000u l=150000u
+  ad=2.73e+11p pd=2.98e+06u as=1.764e+11p ps=1.68e+06u
M1002 a_606_47# a_243_409# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1003 X a_243_409# a_606_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1004 a_243_409# B1 a_225_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.008e+11p ps=1.32e+06u
M1005 a_225_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_243_409# B2 a_137_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A2 a_137_409# VPB phighvt w=1e+06u l=250000u
+  ad=7.95e+11p pd=5.59e+06u as=0p ps=0u
M1008 a_389_47# A1 a_243_409# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_137_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_243_409# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

