* File: sky130_fd_sc_lp__bushold_1.pex.spice
* Created: Wed Sep  2 09:37:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUSHOLD_1%X 1 2 9 15 18 19 22 23 27 28 29 30 31 32
+ 33 34 35 36 48 51
c64 23 0 1.29691e-19 $X=0.65 $Y=1.35
c65 22 0 1.66374e-19 $X=0.65 $Y=1.35
c66 9 0 1.73996e-19 $X=0.715 $Y=0.445
r67 36 68 4.37134 $w=2.88e-07 $l=1.1e-07 $layer=LI1_cond $X=2.17 $Y=2.775
+ $X2=2.17 $Y2=2.885
r68 36 64 9.53746 $w=2.88e-07 $l=2.4e-07 $layer=LI1_cond $X=2.17 $Y=2.775
+ $X2=2.17 $Y2=2.535
r69 35 49 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.45 $X2=2.17
+ $Y2=2.365
r70 35 64 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.45 $X2=2.17
+ $Y2=2.535
r71 35 49 0.914007 $w=2.88e-07 $l=2.3e-08 $layer=LI1_cond $X=2.17 $Y=2.342
+ $X2=2.17 $Y2=2.365
r72 34 35 12.2 $w=2.88e-07 $l=3.07e-07 $layer=LI1_cond $X=2.17 $Y=2.035 $X2=2.17
+ $Y2=2.342
r73 33 34 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=2.035
r74 32 33 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=1.295
+ $X2=2.17 $Y2=1.665
r75 31 32 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=0.925
+ $X2=2.17 $Y2=1.295
r76 30 31 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=0.555
+ $X2=2.17 $Y2=0.925
r77 30 51 4.37134 $w=2.88e-07 $l=1.1e-07 $layer=LI1_cond $X=2.17 $Y=0.555
+ $X2=2.17 $Y2=0.445
r78 28 35 3.3199 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.025 $Y=2.45
+ $X2=2.17 $Y2=2.45
r79 28 29 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=2.025 $Y=2.45
+ $X2=0.815 $Y2=2.45
r80 27 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=2.03
+ $X2=0.65 $Y2=2.195
r81 26 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.65
+ $Y=2.03 $X2=0.65 $Y2=2.03
r82 23 27 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.65 $Y=1.35
+ $X2=0.65 $Y2=2.03
r83 22 26 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.65 $Y=1.35
+ $X2=0.65 $Y2=2.03
r84 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.65
+ $Y=1.35 $X2=0.65 $Y2=1.35
r85 20 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.65 $Y=2.365
+ $X2=0.815 $Y2=2.45
r86 20 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.65 $Y=2.365
+ $X2=0.65 $Y2=2.03
r87 18 19 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=0.762 $Y=2.405
+ $X2=0.762 $Y2=2.555
r88 18 48 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.74 $Y=2.405
+ $X2=0.74 $Y2=2.195
r89 17 23 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.185
+ $X2=0.65 $Y2=1.35
r90 15 19 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.785 $Y=2.885
+ $X2=0.785 $Y2=2.555
r91 9 17 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.715 $Y=0.445
+ $X2=0.715 $Y2=1.185
r92 2 68 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.675 $X2=2.14 $Y2=2.885
r93 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.235 $X2=2.14 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD_1%RESET 3 7 11 12 13 19 22 24
c42 19 0 1.97939e-19 $X=1.19 $Y=1.35
c43 11 0 1.73996e-19 $X=1.2 $Y=1.295
c44 3 0 1.66374e-19 $X=1.145 $Y=0.445
r45 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=2.03
+ $X2=1.19 $Y2=2.195
r46 19 22 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.19 $Y2=2.03
r47 13 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=2.03 $X2=1.19 $Y2=2.03
r48 12 13 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.19 $Y=1.665
+ $X2=1.19 $Y2=2.03
r49 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=1.295
+ $X2=1.19 $Y2=1.665
r50 11 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.35 $X2=1.19 $Y2=1.35
r51 10 19 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.185
+ $X2=1.19 $Y2=1.35
r52 7 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.145 $Y=2.885
+ $X2=1.145 $Y2=2.195
r53 3 10 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.145 $Y=0.445
+ $X2=1.145 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD_1%A_89_535# 1 2 7 9 10 12 14 18 19 20 23 25
+ 29 30 38 40
c72 40 0 3.2763e-19 $X=0.925 $Y=0.84
r73 35 38 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.2 $Y=2.885
+ $X2=0.57 $Y2=2.885
r74 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=2.03 $X2=1.73 $Y2=2.03
r75 30 33 130.408 $w=4.35e-07 $l=1.02e-06 $layer=POLY_cond $X=1.782 $Y=1.01
+ $X2=1.782 $Y2=2.03
r76 29 32 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=1.73 $Y=1.01
+ $X2=1.73 $Y2=2.03
r77 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.01 $X2=1.73 $Y2=1.01
r78 27 29 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=1.73 $Y=0.965
+ $X2=1.73 $Y2=1.01
r79 26 40 5.33677 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=1.055 $Y=0.84
+ $X2=0.925 $Y2=0.84
r80 25 27 6.81649 $w=2.5e-07 $l=1.76777e-07 $layer=LI1_cond $X=1.605 $Y=0.84
+ $X2=1.73 $Y2=0.965
r81 25 26 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=1.605 $Y=0.84
+ $X2=1.055 $Y2=0.84
r82 21 40 1.20171 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=0.925 $Y=0.715
+ $X2=0.925 $Y2=0.84
r83 21 23 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=0.925 $Y=0.715
+ $X2=0.925 $Y2=0.445
r84 19 40 5.33677 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=0.795 $Y=0.84
+ $X2=0.925 $Y2=0.84
r85 19 20 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.795 $Y=0.84
+ $X2=0.315 $Y2=0.84
r86 18 35 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.2 $Y=2.72 $X2=0.2
+ $Y2=2.885
r87 17 20 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=0.2 $Y=0.965
+ $X2=0.315 $Y2=0.84
r88 17 18 87.9364 $w=2.28e-07 $l=1.755e-06 $layer=LI1_cond $X=0.2 $Y=0.965
+ $X2=0.2 $Y2=2.72
r89 16 33 47.9443 $w=4.35e-07 $l=3.75e-07 $layer=POLY_cond $X=1.782 $Y=2.405
+ $X2=1.782 $Y2=2.03
r90 14 30 4.4748 $w=4.35e-07 $l=3.5e-08 $layer=POLY_cond $X=1.782 $Y=0.975
+ $X2=1.782 $Y2=1.01
r91 10 16 27.7985 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.75 $Y=2.655 $X2=1.75
+ $Y2=2.405
r92 10 12 22.172 $w=5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.75 $Y=2.655 $X2=1.75
+ $Y2=2.885
r93 7 14 27.7985 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.75 $Y=0.725 $X2=1.75
+ $Y2=0.975
r94 7 9 26.992 $w=5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.75 $Y=0.725 $X2=1.75
+ $Y2=0.445
r95 2 38 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.445
+ $Y=2.675 $X2=0.57 $Y2=2.885
r96 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.79
+ $Y=0.235 $X2=0.93 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD_1%VPWR 1 6 8 10 17 18 21 27
r26 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.44 $Y2=3.33
r27 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.36 $Y2=3.33
r29 15 17 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.36 $Y2=3.33
r32 10 12 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 8 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.44 $Y2=3.33
r34 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.24
+ $Y2=3.33
r35 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=3.245 $X2=1.36
+ $Y2=3.33
r37 4 6 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.36 $Y=3.245 $X2=1.36
+ $Y2=2.885
r38 1 6 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.675 $X2=1.36 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__BUSHOLD_1%VGND 1 2 9 13 16 17 19 20 21 31 32 38
r33 32 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.44
+ $Y2=0
r34 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 21 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.44
+ $Y2=0
r37 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r38 21 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r39 19 28 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.2
+ $Y2=0
r40 19 20 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.375
+ $Y2=0
r41 18 31 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=2.16
+ $Y2=0
r42 18 20 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.375
+ $Y2=0
r43 16 24 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.335 $Y=0 $X2=0.24
+ $Y2=0
r44 16 17 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.335 $Y=0 $X2=0.48
+ $Y2=0
r45 15 28 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=1.2
+ $Y2=0
r46 15 17 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.48
+ $Y2=0
r47 11 20 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0
r48 11 13 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0.38
r49 7 17 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=0.085
+ $X2=0.48 $Y2=0
r50 7 9 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.48 $Y=0.085
+ $X2=0.48 $Y2=0.38
r51 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.22
+ $Y=0.235 $X2=1.36 $Y2=0.38
r52 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.375
+ $Y=0.235 $X2=0.5 $Y2=0.38
.ends

