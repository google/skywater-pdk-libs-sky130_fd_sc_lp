* File: sky130_fd_sc_lp__a2bb2oi_2.spice
* Created: Wed Sep  2 09:24:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2oi_2.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2oi_2  VNB VPB B1 B2 A1_N A2_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2_N	A2_N
* A1_N	A1_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_B1_M1015_g N_A_113_65#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.8 A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_B2_M1004_g N_A_113_65#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1008 N_Y_M1004_d N_B2_M1008_g N_A_113_65#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.1
+ SB=75004 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_B1_M1018_g N_A_113_65#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=11.424 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_459_39#_M1003_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1 SB=75002.9
+ A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1003_d N_A_459_39#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3717 PD=1.12 PS=1.725 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.5
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1009_s N_A1_N_M1010_g N_A_459_39#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.3717 AS=0.1176 PD=1.725 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.5
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_A1_N_M1019_g N_A_459_39#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1019_d N_A2_N_M1000_g N_A_459_39#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.4
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_A2_N_M1017_g N_A_459_39#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_30_367#_M1002_d N_B1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1005 N_A_30_367#_M1005_d N_B2_M1005_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1012 N_A_30_367#_M1005_d N_B2_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2772 PD=1.54 PS=1.7 NRD=0 NRS=14.0658 M=1 R=8.4 SA=75001.1
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1011 N_A_30_367#_M1011_d N_B1_M1011_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2772 PD=1.54 PS=1.7 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75001.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 N_A_30_367#_M1011_d N_A_459_39#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_A_30_367#_M1016_d N_A_459_39#_M1016_g N_Y_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A1_N_M1001_g N_A_699_367#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1001_d N_A1_N_M1013_g N_A_699_367#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_A_459_39#_M1006_d N_A2_N_M1006_g N_A_699_367#_M1013_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_459_39#_M1006_d N_A2_N_M1014_g N_A_699_367#_M1014_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
c_60 VNB 0 3.08816e-19 $X=0 $Y=0
c_104 VPB 0 1.81764e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a2bb2oi_2.pxi.spice"
*
.ends
*
*
