* File: sky130_fd_sc_lp__and4b_4.pex.spice
* Created: Fri Aug 28 10:08:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4B_4%A_N 3 6 8 9 10 11 12 19 21
r29 19 22 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.707 $Y=1.36
+ $X2=0.707 $Y2=1.525
r30 19 21 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.707 $Y=1.36
+ $X2=0.707 $Y2=1.195
r31 11 12 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=2.035
r32 10 11 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=1.295
+ $X2=0.725 $Y2=1.665
r33 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.36 $X2=0.72 $Y2=1.36
r34 9 10 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=0.925
+ $X2=0.725 $Y2=1.295
r35 8 9 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=0.555
+ $X2=0.725 $Y2=0.925
r36 6 22 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.605 $Y=2.045
+ $X2=0.605 $Y2=1.525
r37 3 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.605 $Y=0.875
+ $X2=0.605 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%A_242_23# 1 2 3 12 16 20 24 28 32 36 40 42
+ 51 53 55 56 60 62 64 66 67 74
c128 66 0 1.19599e-19 $X=2.71 $Y=1.545
c129 40 0 1.95543e-19 $X=2.575 $Y=2.465
r130 71 72 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.715 $Y=1.51
+ $X2=2.145 $Y2=1.51
r131 62 67 16.2203 $w=9.08e-07 $l=4.55e-07 $layer=LI1_cond $X=3.75 $Y=0.71
+ $X2=3.295 $Y2=0.71
r132 62 64 14.144 $w=9.08e-07 $l=1.055e-06 $layer=LI1_cond $X=3.75 $Y=0.71
+ $X2=4.805 $Y2=0.71
r133 58 60 37.7163 $w=3.28e-07 $l=1.08e-06 $layer=LI1_cond $X=3.295 $Y=2.095
+ $X2=4.375 $Y2=2.095
r134 56 58 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.795 $Y=2.095
+ $X2=3.295 $Y2=2.095
r135 55 67 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.795 $Y=1.08
+ $X2=3.295 $Y2=1.08
r136 53 56 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.71 $Y=1.93
+ $X2=2.795 $Y2=2.095
r137 52 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=1.675
+ $X2=2.71 $Y2=1.545
r138 52 53 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.71 $Y=1.675
+ $X2=2.71 $Y2=1.93
r139 51 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=1.415
+ $X2=2.71 $Y2=1.545
r140 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.71 $Y=1.165
+ $X2=2.795 $Y2=1.08
r141 50 51 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.71 $Y=1.165
+ $X2=2.71 $Y2=1.415
r142 49 74 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.52 $Y=1.51
+ $X2=2.575 $Y2=1.51
r143 49 72 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.52 $Y=1.51
+ $X2=2.145 $Y2=1.51
r144 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.51 $X2=2.52 $Y2=1.51
r145 45 71 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.5 $Y=1.51
+ $X2=1.715 $Y2=1.51
r146 45 68 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.5 $Y=1.51
+ $X2=1.285 $Y2=1.51
r147 44 48 45.2112 $w=2.58e-07 $l=1.02e-06 $layer=LI1_cond $X=1.5 $Y=1.545
+ $X2=2.52 $Y2=1.545
r148 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.5
+ $Y=1.51 $X2=1.5 $Y2=1.51
r149 42 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.545
+ $X2=2.71 $Y2=1.545
r150 42 48 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.625 $Y=1.545
+ $X2=2.52 $Y2=1.545
r151 38 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.675
+ $X2=2.575 $Y2=1.51
r152 38 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.575 $Y=1.675
+ $X2=2.575 $Y2=2.465
r153 34 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.345
+ $X2=2.575 $Y2=1.51
r154 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.575 $Y=1.345
+ $X2=2.575 $Y2=0.665
r155 30 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.675
+ $X2=2.145 $Y2=1.51
r156 30 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.145 $Y=1.675
+ $X2=2.145 $Y2=2.465
r157 26 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.345
+ $X2=2.145 $Y2=1.51
r158 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.145 $Y=1.345
+ $X2=2.145 $Y2=0.665
r159 22 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.675
+ $X2=1.715 $Y2=1.51
r160 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.715 $Y=1.675
+ $X2=1.715 $Y2=2.465
r161 18 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.345
+ $X2=1.715 $Y2=1.51
r162 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.715 $Y=1.345
+ $X2=1.715 $Y2=0.665
r163 14 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.675
+ $X2=1.285 $Y2=1.51
r164 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.285 $Y=1.675
+ $X2=1.285 $Y2=2.465
r165 10 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.345
+ $X2=1.285 $Y2=1.51
r166 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.285 $Y=1.345
+ $X2=1.285 $Y2=0.665
r167 3 60 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=1.835 $X2=4.375 $Y2=2.095
r168 2 58 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=1.835 $X2=3.295 $Y2=2.095
r169 1 64 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.665
+ $Y=0.245 $X2=4.805 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%D 3 7 9 12 13
c38 13 0 1.95543e-19 $X=3.06 $Y=1.51
c39 3 0 7.86943e-20 $X=3.08 $Y=2.465
r40 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.51
+ $X2=3.06 $Y2=1.675
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=1.51
+ $X2=3.06 $Y2=1.345
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.51 $X2=3.06 $Y2=1.51
r43 9 13 5.95429 $w=2.98e-07 $l=1.55e-07 $layer=LI1_cond $X=3.115 $Y=1.665
+ $X2=3.115 $Y2=1.51
r44 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.15 $Y=0.665
+ $X2=3.15 $Y2=1.345
r45 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.08 $Y=2.465
+ $X2=3.08 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%C 3 7 9 12 13
c33 13 0 7.86943e-20 $X=3.6 $Y=1.51
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=1.51 $X2=3.6
+ $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=1.51 $X2=3.6
+ $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=1.51 $X2=3.6 $Y2=1.51
r37 9 13 5.3322 $w=3.33e-07 $l=1.55e-07 $layer=LI1_cond $X=3.602 $Y=1.665
+ $X2=3.602 $Y2=1.51
r38 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.51 $Y=2.465
+ $X2=3.51 $Y2=1.675
r39 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.51 $Y=0.665
+ $X2=3.51 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%B 3 7 9 10 14
c34 14 0 1.33412e-19 $X=4.14 $Y=1.51
r35 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.51
+ $X2=4.14 $Y2=1.675
r36 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.51
+ $X2=4.14 $Y2=1.345
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.51 $X2=4.14 $Y2=1.51
r38 10 15 11.6633 $w=4.13e-07 $l=4.2e-07 $layer=LI1_cond $X=4.56 $Y=1.542
+ $X2=4.14 $Y2=1.542
r39 9 15 1.66618 $w=4.13e-07 $l=6e-08 $layer=LI1_cond $X=4.08 $Y=1.542 $X2=4.14
+ $Y2=1.542
r40 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.16 $Y=2.465
+ $X2=4.16 $Y2=1.675
r41 3 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.05 $Y=0.665
+ $X2=4.05 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%A_49_133# 1 2 9 13 16 19 23 24 27 28
c67 27 0 1.33412e-19 $X=4.99 $Y=1.46
r68 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.46 $X2=4.99 $Y2=1.46
r69 25 27 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=4.99 $Y=2.43
+ $X2=4.99 $Y2=1.46
r70 23 25 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.825 $Y=2.52
+ $X2=4.99 $Y2=2.43
r71 23 24 269.263 $w=1.78e-07 $l=4.37e-06 $layer=LI1_cond $X=4.825 $Y=2.52
+ $X2=0.455 $Y2=2.52
r72 19 22 53.9343 $w=2.48e-07 $l=1.17e-06 $layer=LI1_cond $X=0.33 $Y=0.87
+ $X2=0.33 $Y2=2.04
r73 17 24 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=0.33 $Y=2.43
+ $X2=0.455 $Y2=2.52
r74 17 22 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.33 $Y=2.43
+ $X2=0.33 $Y2=2.04
r75 15 28 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=4.665 $Y=1.46
+ $X2=4.99 $Y2=1.46
r76 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.665 $Y=1.46
+ $X2=4.59 $Y2=1.46
r77 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.625
+ $X2=4.59 $Y2=1.46
r78 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.59 $Y=1.625
+ $X2=4.59 $Y2=2.465
r79 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.295
+ $X2=4.59 $Y2=1.46
r80 7 9 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.59 $Y=1.295 $X2=4.59
+ $Y2=0.665
r81 2 22 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.04
r82 1 19 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.665 $X2=0.37 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%VPWR 1 2 3 4 5 18 22 24 28 30 34 38 41 42 43
+ 44 46 47 48 62 63 66 69
r79 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 60 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 60 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r83 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 57 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=3.33
+ $X2=3.725 $Y2=3.33
r85 57 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.89 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 52 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r88 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r89 48 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r90 48 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 48 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 46 59 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.64 $Y=3.33 $X2=4.56
+ $Y2=3.33
r93 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=3.33
+ $X2=4.805 $Y2=3.33
r94 45 62 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.97 $Y=3.33 $X2=5.04
+ $Y2=3.33
r95 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=3.33
+ $X2=4.805 $Y2=3.33
r96 43 55 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.68 $Y2=3.33
r97 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.93 $Y2=3.33
r98 41 51 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.72 $Y2=3.33
r99 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.07 $Y2=3.33
r100 40 55 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=3.33
+ $X2=1.07 $Y2=3.33
r102 36 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.805 $Y=3.245
+ $X2=4.805 $Y2=3.33
r103 36 38 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.805 $Y=3.245
+ $X2=4.805 $Y2=2.9
r104 32 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=3.245
+ $X2=3.725 $Y2=3.33
r105 32 34 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.725 $Y=3.245
+ $X2=3.725 $Y2=2.9
r106 31 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=3.33
+ $X2=2.79 $Y2=3.33
r107 30 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=3.33
+ $X2=3.725 $Y2=3.33
r108 30 31 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.56 $Y=3.33
+ $X2=2.955 $Y2=3.33
r109 26 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=3.33
r110 26 28 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=2.9
r111 25 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.93 $Y2=3.33
r112 24 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.79 $Y2=3.33
r113 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.095 $Y2=3.33
r114 20 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r115 20 22 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.9
r116 16 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r117 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.9
r118 5 38 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=1.835 $X2=4.805 $Y2=2.9
r119 4 34 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.835 $X2=3.725 $Y2=2.9
r120 3 28 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.835 $X2=2.79 $Y2=2.9
r121 2 22 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=2.9
r122 1 18 600 $w=1.7e-07 $l=1.24482e-06 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.835 $X2=1.07 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%X 1 2 3 4 14 15 16 19 21 25 27 28 29 30 37
+ 46
r49 35 37 0.995938 $w=4.03e-07 $l=3.5e-08 $layer=LI1_cond $X=1.165 $Y=2.057
+ $X2=1.2 $Y2=2.057
r50 30 46 5.69108 $w=4.03e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=2.057 $X2=2.36
+ $Y2=2.057
r51 29 30 13.6586 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.057
+ $X2=2.16 $Y2=2.057
r52 29 40 5.12197 $w=4.03e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=2.057
+ $X2=1.5 $Y2=2.057
r53 28 35 2.53308 $w=4.05e-07 $l=9e-08 $layer=LI1_cond $X=1.075 $Y=2.057
+ $X2=1.165 $Y2=2.057
r54 28 40 7.82523 $w=4.03e-07 $l=2.75e-07 $layer=LI1_cond $X=1.225 $Y=2.057
+ $X2=1.5 $Y2=2.057
r55 28 37 0.711385 $w=4.03e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=2.057
+ $X2=1.2 $Y2=2.057
r56 23 25 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.36 $Y=1.075
+ $X2=2.36 $Y2=0.42
r57 22 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.48 $Y2=1.16
r58 21 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.265 $Y=1.16
+ $X2=2.36 $Y2=1.075
r59 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.265 $Y=1.16
+ $X2=1.595 $Y2=1.16
r60 17 27 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.075
+ $X2=1.48 $Y2=1.16
r61 17 19 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.48 $Y=1.075
+ $X2=1.48 $Y2=0.42
r62 15 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.365 $Y=1.16
+ $X2=1.48 $Y2=1.16
r63 15 16 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.365 $Y=1.16
+ $X2=1.165 $Y2=1.16
r64 14 28 5.68537 $w=1.8e-07 $l=2.02e-07 $layer=LI1_cond $X=1.075 $Y=1.855
+ $X2=1.075 $Y2=2.057
r65 13 16 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.075 $Y=1.245
+ $X2=1.165 $Y2=1.16
r66 13 14 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=1.075 $Y=1.245
+ $X2=1.075 $Y2=1.855
r67 4 46 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.835 $X2=2.36 $Y2=2.095
r68 3 40 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.095
r69 2 25 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.22
+ $Y=0.245 $X2=2.36 $Y2=0.42
r70 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.36
+ $Y=0.245 $X2=1.5 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_4%VGND 1 2 3 12 16 20 23 24 26 27 29 30 31 47
+ 48
r63 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r64 45 48 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r65 44 47 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r66 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r67 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r69 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r70 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r71 31 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r72 31 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r73 29 41 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.64
+ $Y2=0
r74 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.865
+ $Y2=0
r75 28 44 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.12
+ $Y2=0
r76 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.865
+ $Y2=0
r77 26 38 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r78 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.93
+ $Y2=0
r79 25 41 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.64
+ $Y2=0
r80 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=1.93
+ $Y2=0
r81 23 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r82 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.09
+ $Y2=0
r83 22 38 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.68
+ $Y2=0
r84 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.09
+ $Y2=0
r85 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0
r86 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0.37
r87 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0
r88 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.93 $Y=0.085
+ $X2=1.93 $Y2=0.39
r89 10 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=0.085
+ $X2=1.09 $Y2=0
r90 10 12 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=1.09 $Y=0.085
+ $X2=1.09 $Y2=0.39
r91 3 20 91 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=2 $X=2.65
+ $Y=0.245 $X2=2.865 $Y2=0.37
r92 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.79
+ $Y=0.245 $X2=1.93 $Y2=0.39
r93 1 12 91 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=2 $X=0.68
+ $Y=0.665 $X2=1.07 $Y2=0.39
.ends

