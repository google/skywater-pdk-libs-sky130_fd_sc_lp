* File: sky130_fd_sc_lp__busreceiver_m.pex.spice
* Created: Wed Sep  2 09:38:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_M%A_47_178# 1 2 8 9 11 14 18 20 23 27 30
+ 32 35
r57 36 38 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.31 $Y=2.015
+ $X2=0.475 $Y2=2.015
r58 32 34 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=0.495
+ $X2=1.12 $Y2=0.66
r59 30 35 4.70473 $w=1.9e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.14 $Y=1.93
+ $X2=1.12 $Y2=2.015
r60 30 34 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=1.14 $Y=1.93
+ $X2=1.14 $Y2=0.66
r61 25 35 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.1 $X2=1.12
+ $Y2=2.015
r62 25 27 36.7056 $w=2.08e-07 $l=6.95e-07 $layer=LI1_cond $X=1.12 $Y=2.1
+ $X2=1.12 $Y2=2.795
r63 23 38 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.71 $Y=2.015
+ $X2=0.475 $Y2=2.015
r64 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=2.015 $X2=0.71 $Y2=2.015
r65 20 35 1.74598 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.015 $Y=2.015
+ $X2=1.12 $Y2=2.015
r66 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.015 $Y=2.015
+ $X2=0.71 $Y2=2.015
r67 16 18 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.31 $Y=0.965
+ $X2=0.475 $Y2=0.965
r68 12 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.18
+ $X2=0.475 $Y2=2.015
r69 12 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.475 $Y=2.18
+ $X2=0.475 $Y2=2.86
r70 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=0.89
+ $X2=0.475 $Y2=0.965
r71 9 11 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.475 $Y=0.89
+ $X2=0.475 $Y2=0.56
r72 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.31 $Y=1.85
+ $X2=0.31 $Y2=2.015
r73 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.04 $X2=0.31
+ $Y2=0.965
r74 7 8 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.31 $Y=1.04 $X2=0.31
+ $Y2=1.85
r75 2 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.65 $X2=1.12 $Y2=2.795
r76 1 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.35 $X2=1.12 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_M%A 3 5 7 9 12 14 15 16 25
r46 24 25 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=0.905 $Y=1.445
+ $X2=1.19 $Y2=1.445
r47 21 24 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=0.79 $Y=1.445
+ $X2=0.905 $Y2=1.445
r48 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.79
+ $Y=1.445 $X2=0.79 $Y2=1.445
r49 16 22 10.5641 $w=2.38e-07 $l=2.2e-07 $layer=LI1_cond $X=0.755 $Y=1.665
+ $X2=0.755 $Y2=1.445
r50 15 22 7.20277 $w=2.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.755 $Y=1.295
+ $X2=0.755 $Y2=1.445
r51 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=0.925
+ $X2=0.755 $Y2=1.295
r52 10 12 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.905 $Y=2.465
+ $X2=1.19 $Y2=2.465
r53 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.19 $Y=2.39 $X2=1.19
+ $Y2=2.465
r54 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.61
+ $X2=1.19 $Y2=1.445
r55 8 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.19 $Y=1.61 $X2=1.19
+ $Y2=2.39
r56 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=2.54
+ $X2=0.905 $Y2=2.465
r57 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=2.54
+ $X2=0.905 $Y2=2.86
r58 1 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.28
+ $X2=0.905 $Y2=1.445
r59 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.905 $Y=1.28
+ $X2=0.905 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_M%X 1 2 7 8 9 10 11 12 20
r16 11 12 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r17 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.035
+ $X2=0.26 $Y2=2.405
r18 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r19 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295 $X2=0.26
+ $Y2=1.665
r20 7 8 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.925 $X2=0.26
+ $Y2=1.295
r21 7 20 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=0.26 $Y=0.925 $X2=0.26
+ $Y2=0.625
r22 2 12 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.65 $X2=0.26 $Y2=2.795
r23 1 20 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.35 $X2=0.26 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_M%VPWR 1 6 9 10 11 18 19
r19 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r20 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r22 11 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 9 14 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 9 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.69 $Y2=3.33
r25 8 18 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=1.2 $Y2=3.33
r26 8 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.69 $Y2=3.33
r27 4 10 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r28 4 6 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.925
r29 1 6 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.65 $X2=0.69 $Y2=2.925
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_M%VGND 1 6 9 10 11 18 19
r19 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r20 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r21 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r22 11 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r23 9 14 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r24 9 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.69
+ $Y2=0
r25 8 18 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r26 8 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.69
+ $Y2=0
r27 4 10 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r28 4 6 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0.495
r29 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.35 $X2=0.69 $Y2=0.495
.ends

