* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_273_49# B2 a_179_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_549_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_96_49# C1 a_179_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_287_367# B2 a_96_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_96_49# A2 a_549_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A2 a_273_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_273_49# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR B1 a_287_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_179_49# B1 a_273_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND a_96_49# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_96_49# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR a_96_49# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
