* File: sky130_fd_sc_lp__o32a_2.spice
* Created: Fri Aug 28 11:17:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32a_2.pex.spice"
.subckt sky130_fd_sc_lp__o32a_2  VNB VPB A1 A2 A3 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_85_21#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_85_21#_M1013_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.231 AS=0.1176 PD=1.39 PS=1.12 NRD=18.564 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1001 N_A_341_47#_M1001_d N_A1_M1001_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.231 PD=1.12 PS=1.39 NRD=0 NRS=19.992 M=1 R=5.6 SA=75001.3
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_341_47#_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=1.41 PS=1.12 NRD=19.992 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1003 N_A_341_47#_M1003_d N_A3_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=1.41 NRD=0 NRS=21.42 M=1 R=5.6 SA=75002.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_A_85_21#_M1009_d N_B2_M1009_g N_A_341_47#_M1003_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6
+ SA=75002.9 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1007 N_A_341_47#_M1007_d N_B1_M1007_g N_A_85_21#_M1009_d VNB NSHORT L=0.15
+ W=0.84 AD=0.252 AS=0.1344 PD=2.28 PS=1.16 NRD=2.136 NRS=0 M=1 R=5.6 SA=75003.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_X_M1006_d N_A_85_21#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1012 N_X_M1006_d N_A_85_21#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1000 A_355_367# N_A1_M1000_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3906 PD=1.47 PS=1.88 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1008 A_427_367# N_A2_M1008_g A_355_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75001.8
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1005 N_A_85_21#_M1005_d N_A3_M1005_g A_427_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=7.8012 NRS=21.8867 M=1 R=8.4
+ SA=75002.3 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1010 A_643_367# N_B2_M1010_g N_A_85_21#_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=9.3772 M=1 R=8.4
+ SA=75002.8 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g A_643_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75003.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o32a_2.pxi.spice"
*
.ends
*
*
