* File: sky130_fd_sc_lp__sdfrbp_1.spice
* Created: Fri Aug 28 11:27:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrbp_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfrbp_1  VNB VPB SCE D SCD CLK RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1042 N_VGND_M1042_d N_SCE_M1042_g N_A_27_75#_M1042_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 noxref_26 N_A_27_75#_M1029_g N_noxref_25_M1029_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.1113 PD=0.81 PS=1.37 NRD=37.14 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_367_491#_M1011_d N_D_M1011_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0777 PD=0.7 PS=0.81 NRD=0 NRS=37.14 M=1 R=2.8 SA=75000.7
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1038 noxref_27 N_SCE_M1038_g N_A_367_491#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1030 N_noxref_25_M1030_d N_SCD_M1030_g noxref_27 VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_RESET_B_M1021_g N_noxref_25_M1030_d VNB NSHORT L=0.15
+ W=0.42 AD=0.2145 AS=0.0735 PD=1.36 PS=0.77 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1021_d N_CLK_M1015_g N_A_840_119#_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.2145 AS=0.0588 PD=1.36 PS=0.7 NRD=130.2 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_840_119#_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.103375 AS=0.0588 PD=0.975 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_1024_367#_M1013_d N_A_840_119#_M1013_g N_VGND_M1023_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.103375 PD=0.7 PS=0.975 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75002.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_1024_367#_M1013_d N_A_840_119#_M1018_g N_VGND_M1018_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1239 PD=0.7 PS=1.43 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_A_1246_463#_M1031_d N_A_840_119#_M1031_g N_A_367_491#_M1031_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1033 A_1430_119# N_A_1024_367#_M1033_g N_A_1246_463#_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1026 A_1502_119# N_A_1374_362#_M1026_g A_1430_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_RESET_B_M1014_g A_1502_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.127783 AS=0.0441 PD=0.939057 PS=0.63 NRD=71.208 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_1374_362#_M1004_d N_A_1246_463#_M1004_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2289 AS=0.194717 PD=1.51 PS=1.43094 NRD=56.748 NRS=23.436
+ M=1 R=4.26667 SA=75001.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1043 N_A_1812_379#_M1043_d N_A_1024_367#_M1043_g N_A_1374_362#_M1004_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.144604 AS=0.2289 PD=1.25585 PS=1.51 NRD=22.488
+ NRS=56.748 M=1 R=4.26667 SA=75002.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1024 A_1960_68# N_A_840_119#_M1024_g N_A_1812_379#_M1043_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0948962 PD=0.63 PS=0.824151 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_2002_42#_M1019_g A_1960_68# VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0441 PD=0.8 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1027 A_2138_68# N_RESET_B_M1027_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0798 PD=0.63 PS=0.8 NRD=14.28 NRS=28.56 M=1 R=2.8 SA=75003.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_2002_42#_M1005_d N_A_1812_379#_M1005_g A_2138_68# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1036 N_A_2352_327#_M1036_d N_A_1812_379#_M1036_g N_VGND_M1036_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_2352_327#_M1008_g N_Q_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1034 N_Q_N_M1034_d N_A_1812_379#_M1034_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_SCE_M1000_g N_A_27_75#_M1000_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1020 A_295_491# N_SCE_M1020_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1028 N_A_367_491#_M1028_d N_D_M1028_g A_295_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1009 A_453_491# N_A_27_75#_M1009_g N_A_367_491#_M1028_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1104 AS=0.0896 PD=0.985 PS=0.92 NRD=36.1495 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_VPWR_M1017_d N_SCD_M1017_g A_453_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.1104 PD=1.03 PS=0.985 NRD=12.2928 NRS=36.1495 M=1 R=4.26667
+ SA=75001.9 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1040 N_A_367_491#_M1040_d N_RESET_B_M1040_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=21.5321 M=1 R=4.26667
+ SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_CLK_M1001_g N_A_840_119#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_A_1024_367#_M1006_d N_A_840_119#_M1006_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1022 N_A_1246_463#_M1022_d N_A_1024_367#_M1022_g N_A_367_491#_M1022_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1449 PD=0.7 PS=1.53 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.3 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 A_1332_463# N_A_840_119#_M1007_g N_A_1246_463#_M1022_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1037 N_VPWR_M1037_d N_A_1374_362#_M1037_g A_1332_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1332 AS=0.0441 PD=1.11 PS=0.63 NRD=39.8531 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_1246_463#_M1010_d N_RESET_B_M1010_g N_VPWR_M1037_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1332 PD=1.37 PS=1.11 NRD=0 NRS=122.948 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_1374_362#_M1012_d N_A_1246_463#_M1012_g N_VPWR_M1012_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1041 N_A_1812_379#_M1041_d N_A_840_119#_M1041_g N_A_1374_362#_M1012_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2419 AS=0.1176 PD=2.08 PS=1.12 NRD=37.5088 NRS=0
+ M=1 R=5.6 SA=75000.6 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1003 A_1953_496# N_A_1024_367#_M1003_g N_A_1812_379#_M1041_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.08505 AS=0.12095 PD=0.825 PS=1.04 NRD=69.1667 NRS=56.2829
+ M=1 R=2.8 SA=75001 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_2002_42#_M1032_g A_1953_496# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0739375 AS=0.08505 PD=0.81 PS=0.825 NRD=9.3772 NRS=69.1667 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1002 N_A_2002_42#_M1002_d N_RESET_B_M1002_g N_VPWR_M1032_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0739375 PD=0.7 PS=0.81 NRD=0 NRS=11.7215 M=1 R=2.8
+ SA=75001.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_1812_379#_M1025_g N_A_2002_42#_M1002_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.126 AS=0.0588 PD=1.44 PS=0.7 NRD=16.4101 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_A_2352_327#_M1035_d N_A_1812_379#_M1035_g N_VPWR_M1035_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1984 PD=1.81 PS=1.9 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1039 N_VPWR_M1039_d N_A_2352_327#_M1039_g N_Q_M1039_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_Q_N_M1016_d N_A_1812_379#_M1016_g N_VPWR_M1039_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX44_noxref VNB VPB NWDIODE A=26.8865 P=32.73
c_2054 A_1332_463# 0 3.01024e-19 $X=6.66 $Y=2.315
*
.include "sky130_fd_sc_lp__sdfrbp_1.pxi.spice"
*
.ends
*
*
