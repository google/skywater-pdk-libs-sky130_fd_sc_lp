* File: sky130_fd_sc_lp__and4b_1.pxi.spice
* Created: Wed Sep  2 09:33:27 2020
* 
x_PM_SKY130_FD_SC_LP__AND4B_1%A_N N_A_N_M1005_g N_A_N_M1010_g N_A_N_c_87_n
+ N_A_N_c_88_n A_N N_A_N_c_89_n N_A_N_c_90_n PM_SKY130_FD_SC_LP__AND4B_1%A_N
x_PM_SKY130_FD_SC_LP__AND4B_1%A_27_49# N_A_27_49#_M1005_s N_A_27_49#_M1010_s
+ N_A_27_49#_M1008_g N_A_27_49#_c_119_n N_A_27_49#_c_120_n N_A_27_49#_c_121_n
+ N_A_27_49#_M1001_g N_A_27_49#_c_122_n N_A_27_49#_c_123_n N_A_27_49#_c_131_n
+ N_A_27_49#_c_124_n N_A_27_49#_c_125_n N_A_27_49#_c_132_n N_A_27_49#_c_133_n
+ N_A_27_49#_c_126_n N_A_27_49#_c_127_n N_A_27_49#_c_128_n N_A_27_49#_c_129_n
+ PM_SKY130_FD_SC_LP__AND4B_1%A_27_49#
x_PM_SKY130_FD_SC_LP__AND4B_1%B N_B_M1002_g N_B_M1003_g B B N_B_c_202_n
+ PM_SKY130_FD_SC_LP__AND4B_1%B
x_PM_SKY130_FD_SC_LP__AND4B_1%C N_C_M1004_g N_C_M1009_g C C N_C_c_238_n
+ PM_SKY130_FD_SC_LP__AND4B_1%C
x_PM_SKY130_FD_SC_LP__AND4B_1%D N_D_c_273_n N_D_M1011_g N_D_M1007_g D D
+ N_D_c_278_n PM_SKY130_FD_SC_LP__AND4B_1%D
x_PM_SKY130_FD_SC_LP__AND4B_1%A_215_367# N_A_215_367#_M1001_s
+ N_A_215_367#_M1008_d N_A_215_367#_M1009_d N_A_215_367#_M1006_g
+ N_A_215_367#_M1000_g N_A_215_367#_c_317_n N_A_215_367#_c_318_n
+ N_A_215_367#_c_319_n N_A_215_367#_c_320_n N_A_215_367#_c_321_n
+ N_A_215_367#_c_322_n N_A_215_367#_c_323_n N_A_215_367#_c_324_n
+ N_A_215_367#_c_331_n N_A_215_367#_c_325_n N_A_215_367#_c_326_n
+ N_A_215_367#_c_327_n PM_SKY130_FD_SC_LP__AND4B_1%A_215_367#
x_PM_SKY130_FD_SC_LP__AND4B_1%VPWR N_VPWR_M1010_d N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n VPWR
+ N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_416_n
+ N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n PM_SKY130_FD_SC_LP__AND4B_1%VPWR
x_PM_SKY130_FD_SC_LP__AND4B_1%X N_X_M1006_d N_X_M1000_d X X X X X X X
+ N_X_c_464_n X PM_SKY130_FD_SC_LP__AND4B_1%X
x_PM_SKY130_FD_SC_LP__AND4B_1%VGND N_VGND_M1005_d N_VGND_M1011_d N_VGND_c_482_n
+ N_VGND_c_483_n VGND N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n
+ N_VGND_c_487_n N_VGND_c_488_n PM_SKY130_FD_SC_LP__AND4B_1%VGND
cc_1 VNB N_A_N_M1005_g 0.0339975f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_2 VNB N_A_N_M1010_g 0.00491479f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.045
cc_3 VNB N_A_N_c_87_n 0.0269388f $X=-0.19 $Y=-0.245 $X2=0.412 $Y2=1.445
cc_4 VNB N_A_N_c_88_n 0.0233151f $X=-0.19 $Y=-0.245 $X2=0.412 $Y2=1.595
cc_5 VNB N_A_N_c_89_n 0.0194255f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_6 VNB N_A_N_c_90_n 0.0235866f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_7 VNB N_A_27_49#_M1008_g 0.0103948f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_8 VNB N_A_27_49#_c_119_n 0.0220998f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.445
cc_9 VNB N_A_27_49#_c_120_n 0.0165034f $X=-0.19 $Y=-0.245 $X2=0.412 $Y2=1.445
cc_10 VNB N_A_27_49#_c_121_n 0.019435f $X=-0.19 $Y=-0.245 $X2=0.412 $Y2=1.595
cc_11 VNB N_A_27_49#_c_122_n 0.0166813f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_12 VNB N_A_27_49#_c_123_n 0.0140007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_49#_c_124_n 0.0101958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_49#_c_125_n 0.0114438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_49#_c_126_n 0.00379819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_49#_c_127_n 0.0258184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_49#_c_128_n 0.0017728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_49#_c_129_n 0.00100303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_M1002_g 0.00640127f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_20 VNB N_B_M1003_g 0.0379742f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.045
cc_21 VNB B 0.0026628f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_22 VNB N_B_c_202_n 0.04683f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_23 VNB N_C_M1004_g 0.0415362f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_24 VNB C 0.00519658f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_25 VNB N_C_c_238_n 0.0287159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_D_c_273_n 0.0410926f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.925
cc_27 VNB N_D_M1011_g 0.0287286f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_28 VNB N_D_M1007_g 0.0163261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_215_367#_M1000_g 0.00834375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_215_367#_c_317_n 0.00268544f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_31 VNB N_A_215_367#_c_318_n 0.00303734f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_32 VNB N_A_215_367#_c_319_n 0.00585758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_215_367#_c_320_n 0.0220576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_215_367#_c_321_n 8.26067e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_215_367#_c_322_n 0.0010459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_215_367#_c_323_n 0.00538903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_215_367#_c_324_n 0.0333424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_215_367#_c_325_n 0.00184091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_215_367#_c_326_n 0.00219462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_215_367#_c_327_n 0.0214511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_416_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB X 0.00826307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB X 0.0325046f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_44 VNB N_X_c_464_n 0.0243299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_482_n 0.00560572f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_46 VNB N_VGND_c_483_n 0.00442308f $X=-0.19 $Y=-0.245 $X2=0.412 $Y2=1.595
cc_47 VNB N_VGND_c_484_n 0.0148678f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.09
cc_48 VNB N_VGND_c_485_n 0.0631519f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.26
cc_49 VNB N_VGND_c_486_n 0.0190369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_487_n 0.211165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_488_n 0.00517829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_A_N_M1010_g 0.029773f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.045
cc_53 VPB N_A_27_49#_M1008_g 0.0234501f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.09
cc_54 VPB N_A_27_49#_c_131_n 0.0145966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_27_49#_c_132_n 0.00543328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_27_49#_c_133_n 0.0095003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_27_49#_c_128_n 3.70661e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B_M1002_g 0.0267031f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.455
cc_59 VPB B 0.00478812f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.09
cc_60 VPB N_C_M1009_g 0.0262867f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.045
cc_61 VPB C 0.00327157f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.09
cc_62 VPB N_C_c_238_n 0.00924845f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_D_M1007_g 0.0320992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB D 0.00772763f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.445
cc_65 VPB N_D_c_278_n 0.0484203f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.26
cc_66 VPB N_A_215_367#_M1000_g 0.0258113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_215_367#_c_319_n 0.00135015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_215_367#_c_322_n 0.0015979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_215_367#_c_331_n 0.00447255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_417_n 0.048323f $X=-0.19 $Y=1.655 $X2=0.412 $Y2=1.445
cc_71 VPB N_VPWR_c_418_n 0.044377f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.09
cc_72 VPB N_VPWR_c_419_n 0.00940087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_420_n 0.00369332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_421_n 0.0212365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_422_n 0.0207798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_423_n 0.0177201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_424_n 0.0164025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_416_n 0.105875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_426_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_427_n 0.0141117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_428_n 0.00497525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB X 0.0087145f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.09
cc_83 VPB X 0.00955129f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.445
cc_84 VPB X 0.0450697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 N_A_N_c_88_n N_A_27_49#_M1008_g 0.0222421f $X=0.412 $Y=1.595 $X2=0 $Y2=0
cc_86 N_A_N_M1005_g N_A_27_49#_c_120_n 0.0106296f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_87 N_A_N_c_87_n N_A_27_49#_c_122_n 0.0106296f $X=0.412 $Y=1.445 $X2=0 $Y2=0
cc_88 N_A_N_M1005_g N_A_27_49#_c_124_n 0.0143664f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_89 N_A_N_c_88_n N_A_27_49#_c_124_n 0.00143229f $X=0.412 $Y=1.595 $X2=0 $Y2=0
cc_90 N_A_N_c_89_n N_A_27_49#_c_124_n 0.0012716f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_91 N_A_N_c_90_n N_A_27_49#_c_124_n 0.013916f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_92 N_A_N_c_89_n N_A_27_49#_c_125_n 0.0039342f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_93 N_A_N_c_90_n N_A_27_49#_c_125_n 0.0166219f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_94 N_A_N_M1010_g N_A_27_49#_c_132_n 0.017247f $X=0.53 $Y=2.045 $X2=0 $Y2=0
cc_95 N_A_N_c_88_n N_A_27_49#_c_132_n 7.15875e-19 $X=0.412 $Y=1.595 $X2=0 $Y2=0
cc_96 N_A_N_c_90_n N_A_27_49#_c_132_n 0.00853968f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_97 N_A_N_c_88_n N_A_27_49#_c_133_n 0.00612622f $X=0.412 $Y=1.595 $X2=0 $Y2=0
cc_98 N_A_N_c_90_n N_A_27_49#_c_133_n 0.022679f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_99 N_A_N_M1005_g N_A_27_49#_c_126_n 0.00399646f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_100 N_A_N_c_89_n N_A_27_49#_c_126_n 7.84456e-19 $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_101 N_A_N_c_90_n N_A_27_49#_c_126_n 0.0343531f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_102 N_A_N_c_89_n N_A_27_49#_c_127_n 0.0106296f $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_103 N_A_N_c_90_n N_A_27_49#_c_127_n 5.11391e-19 $X=0.385 $Y=1.09 $X2=0 $Y2=0
cc_104 N_A_N_c_88_n N_A_27_49#_c_128_n 0.00446112f $X=0.412 $Y=1.595 $X2=0 $Y2=0
cc_105 N_A_N_c_87_n N_A_27_49#_c_129_n 7.84456e-19 $X=0.412 $Y=1.445 $X2=0 $Y2=0
cc_106 N_A_N_M1005_g N_A_215_367#_c_318_n 0.00290041f $X=0.475 $Y=0.455 $X2=0
+ $Y2=0
cc_107 N_A_N_M1010_g N_VPWR_c_417_n 0.0106119f $X=0.53 $Y=2.045 $X2=0 $Y2=0
cc_108 N_A_N_M1005_g N_VGND_c_482_n 0.0102049f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_109 N_A_N_M1005_g N_VGND_c_484_n 0.00348975f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_110 N_A_N_M1005_g N_VGND_c_487_n 0.00511446f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_111 N_A_27_49#_c_121_n N_B_M1003_g 0.0503454f $X=1.425 $Y=0.775 $X2=0 $Y2=0
cc_112 N_A_27_49#_c_127_n N_B_M1003_g 0.00390192f $X=0.98 $Y=0.94 $X2=0 $Y2=0
cc_113 N_A_27_49#_M1008_g N_B_c_202_n 0.0253373f $X=1 $Y=2.045 $X2=0 $Y2=0
cc_114 N_A_27_49#_c_119_n N_B_c_202_n 0.00650162f $X=1.35 $Y=0.85 $X2=0 $Y2=0
cc_115 N_A_27_49#_c_126_n N_B_c_202_n 2.03482e-19 $X=0.98 $Y=0.94 $X2=0 $Y2=0
cc_116 N_A_27_49#_c_127_n N_B_c_202_n 0.0145502f $X=0.98 $Y=0.94 $X2=0 $Y2=0
cc_117 N_A_27_49#_c_128_n N_B_c_202_n 2.21826e-19 $X=0.845 $Y=1.695 $X2=0 $Y2=0
cc_118 N_A_27_49#_c_119_n N_A_215_367#_c_317_n 4.0101e-19 $X=1.35 $Y=0.85 $X2=0
+ $Y2=0
cc_119 N_A_27_49#_c_120_n N_A_215_367#_c_317_n 0.00591521f $X=1.145 $Y=0.85
+ $X2=0 $Y2=0
cc_120 N_A_27_49#_c_121_n N_A_215_367#_c_317_n 0.00531989f $X=1.425 $Y=0.775
+ $X2=0 $Y2=0
cc_121 N_A_27_49#_c_124_n N_A_215_367#_c_317_n 0.00163502f $X=0.76 $Y=0.74 $X2=0
+ $Y2=0
cc_122 N_A_27_49#_c_119_n N_A_215_367#_c_318_n 0.00560126f $X=1.35 $Y=0.85 $X2=0
+ $Y2=0
cc_123 N_A_27_49#_c_121_n N_A_215_367#_c_318_n 0.00854668f $X=1.425 $Y=0.775
+ $X2=0 $Y2=0
cc_124 N_A_27_49#_c_124_n N_A_215_367#_c_318_n 0.0144356f $X=0.76 $Y=0.74 $X2=0
+ $Y2=0
cc_125 N_A_27_49#_c_126_n N_A_215_367#_c_318_n 0.00250451f $X=0.98 $Y=0.94 $X2=0
+ $Y2=0
cc_126 N_A_27_49#_M1008_g N_A_215_367#_c_319_n 0.002515f $X=1 $Y=2.045 $X2=0
+ $Y2=0
cc_127 N_A_27_49#_c_132_n N_A_215_367#_c_319_n 0.00514526f $X=0.76 $Y=1.78 $X2=0
+ $Y2=0
cc_128 N_A_27_49#_c_126_n N_A_215_367#_c_319_n 0.0308883f $X=0.98 $Y=0.94 $X2=0
+ $Y2=0
cc_129 N_A_27_49#_c_127_n N_A_215_367#_c_319_n 0.00343494f $X=0.98 $Y=0.94 $X2=0
+ $Y2=0
cc_130 N_A_27_49#_c_128_n N_A_215_367#_c_319_n 0.0115305f $X=0.845 $Y=1.695
+ $X2=0 $Y2=0
cc_131 N_A_27_49#_M1008_g N_A_215_367#_c_331_n 3.02405e-19 $X=1 $Y=2.045 $X2=0
+ $Y2=0
cc_132 N_A_27_49#_c_122_n N_A_215_367#_c_331_n 0.00127086f $X=0.98 $Y=1.445
+ $X2=0 $Y2=0
cc_133 N_A_27_49#_c_132_n N_A_215_367#_c_331_n 0.00429429f $X=0.76 $Y=1.78 $X2=0
+ $Y2=0
cc_134 N_A_27_49#_c_119_n N_A_215_367#_c_325_n 0.00721496f $X=1.35 $Y=0.85 $X2=0
+ $Y2=0
cc_135 N_A_27_49#_c_126_n N_A_215_367#_c_325_n 0.0139285f $X=0.98 $Y=0.94 $X2=0
+ $Y2=0
cc_136 N_A_27_49#_c_127_n N_A_215_367#_c_325_n 0.00125597f $X=0.98 $Y=0.94 $X2=0
+ $Y2=0
cc_137 N_A_27_49#_c_132_n N_VPWR_M1010_d 0.00222628f $X=0.76 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_27_49#_M1008_g N_VPWR_c_417_n 0.00717747f $X=1 $Y=2.045 $X2=0 $Y2=0
cc_139 N_A_27_49#_c_122_n N_VPWR_c_417_n 2.87063e-19 $X=0.98 $Y=1.445 $X2=0
+ $Y2=0
cc_140 N_A_27_49#_c_132_n N_VPWR_c_417_n 0.018233f $X=0.76 $Y=1.78 $X2=0 $Y2=0
cc_141 N_A_27_49#_c_124_n N_VGND_M1005_d 0.00214584f $X=0.76 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_27_49#_c_120_n N_VGND_c_482_n 2.22223e-19 $X=1.145 $Y=0.85 $X2=0
+ $Y2=0
cc_143 N_A_27_49#_c_121_n N_VGND_c_482_n 0.00231444f $X=1.425 $Y=0.775 $X2=0
+ $Y2=0
cc_144 N_A_27_49#_c_124_n N_VGND_c_482_n 0.0214787f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_27_49#_c_123_n N_VGND_c_484_n 0.0142975f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_146 N_A_27_49#_c_124_n N_VGND_c_484_n 0.00235807f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_27_49#_c_120_n N_VGND_c_485_n 5.87535e-19 $X=1.145 $Y=0.85 $X2=0
+ $Y2=0
cc_148 N_A_27_49#_c_121_n N_VGND_c_485_n 0.00357877f $X=1.425 $Y=0.775 $X2=0
+ $Y2=0
cc_149 N_A_27_49#_c_124_n N_VGND_c_485_n 0.00368443f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_27_49#_M1005_s N_VGND_c_487_n 0.00231058f $X=0.135 $Y=0.245 $X2=0
+ $Y2=0
cc_151 N_A_27_49#_c_121_n N_VGND_c_487_n 0.00648295f $X=1.425 $Y=0.775 $X2=0
+ $Y2=0
cc_152 N_A_27_49#_c_123_n N_VGND_c_487_n 0.00978901f $X=0.26 $Y=0.455 $X2=0
+ $Y2=0
cc_153 N_A_27_49#_c_124_n N_VGND_c_487_n 0.0114233f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_154 N_B_M1003_g N_C_M1004_g 0.0456269f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_155 B N_C_M1004_g 3.82374e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 B N_C_M1009_g 3.06317e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_157 N_B_M1003_g C 0.00203794f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_158 B C 0.0439217f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_B_M1002_g N_C_c_238_n 0.0020338f $X=1.43 $Y=2.045 $X2=0 $Y2=0
cc_160 B N_C_c_238_n 5.65594e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B_c_202_n N_C_c_238_n 0.0456269f $X=1.785 $Y=1.375 $X2=0 $Y2=0
cc_162 N_B_M1003_g N_A_215_367#_c_318_n 0.00476187f $X=1.785 $Y=0.445 $X2=0
+ $Y2=0
cc_163 N_B_M1002_g N_A_215_367#_c_319_n 0.00601515f $X=1.43 $Y=2.045 $X2=0 $Y2=0
cc_164 N_B_M1003_g N_A_215_367#_c_319_n 0.00344014f $X=1.785 $Y=0.445 $X2=0
+ $Y2=0
cc_165 B N_A_215_367#_c_319_n 0.0400387f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B_c_202_n N_A_215_367#_c_319_n 0.00829296f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_167 N_B_M1003_g N_A_215_367#_c_320_n 0.0120457f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_168 B N_A_215_367#_c_320_n 0.0207452f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B_c_202_n N_A_215_367#_c_320_n 0.00318273f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_170 N_B_M1002_g N_A_215_367#_c_331_n 0.0112086f $X=1.43 $Y=2.045 $X2=0 $Y2=0
cc_171 N_B_c_202_n N_A_215_367#_c_325_n 0.00324503f $X=1.785 $Y=1.375 $X2=0
+ $Y2=0
cc_172 N_B_M1002_g N_VPWR_c_417_n 7.10841e-19 $X=1.43 $Y=2.045 $X2=0 $Y2=0
cc_173 N_B_M1002_g N_VPWR_c_418_n 0.0121231f $X=1.43 $Y=2.045 $X2=0 $Y2=0
cc_174 B N_VPWR_c_418_n 0.0247121f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_175 N_B_c_202_n N_VPWR_c_418_n 0.00129012f $X=1.785 $Y=1.375 $X2=0 $Y2=0
cc_176 N_B_M1003_g N_VGND_c_485_n 0.00585385f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_177 N_B_M1003_g N_VGND_c_487_n 0.00624738f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_178 N_C_M1004_g N_D_c_273_n 0.00479939f $X=2.145 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_179 C N_D_c_273_n 2.66765e-19 $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_180 N_C_c_238_n N_D_c_273_n 5.45698e-19 $X=2.235 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_181 N_C_M1004_g N_D_M1011_g 0.064383f $X=2.145 $Y=0.445 $X2=0 $Y2=0
cc_182 N_C_M1004_g N_D_M1007_g 8.30702e-19 $X=2.145 $Y=0.445 $X2=0 $Y2=0
cc_183 C N_D_M1007_g 4.29063e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_184 N_C_c_238_n N_D_M1007_g 0.0282668f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_185 N_C_M1009_g D 6.74439e-19 $X=2.37 $Y=2.045 $X2=0 $Y2=0
cc_186 C N_A_215_367#_c_319_n 3.13535e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_187 N_C_M1004_g N_A_215_367#_c_320_n 0.0110984f $X=2.145 $Y=0.445 $X2=0 $Y2=0
cc_188 C N_A_215_367#_c_320_n 0.0227288f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_189 N_C_c_238_n N_A_215_367#_c_320_n 0.00433001f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_190 N_C_M1004_g N_A_215_367#_c_321_n 0.0019957f $X=2.145 $Y=0.445 $X2=0 $Y2=0
cc_191 C N_A_215_367#_c_322_n 0.019032f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_192 N_C_c_238_n N_A_215_367#_c_322_n 0.00378997f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_193 N_C_M1004_g N_A_215_367#_c_326_n 8.95814e-19 $X=2.145 $Y=0.445 $X2=0
+ $Y2=0
cc_194 C N_A_215_367#_c_326_n 0.0269171f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_195 N_C_c_238_n N_A_215_367#_c_326_n 0.00151988f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_196 N_C_M1009_g N_VPWR_c_418_n 0.0104502f $X=2.37 $Y=2.045 $X2=0 $Y2=0
cc_197 C N_VPWR_c_418_n 0.023321f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_198 N_C_c_238_n N_VPWR_c_418_n 0.0013052f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_199 N_C_M1004_g N_VGND_c_485_n 0.00890921f $X=2.145 $Y=0.445 $X2=0 $Y2=0
cc_200 N_C_M1004_g N_VGND_c_487_n 0.00624738f $X=2.145 $Y=0.445 $X2=0 $Y2=0
cc_201 N_D_M1007_g N_A_215_367#_M1000_g 0.0217856f $X=2.8 $Y=2.045 $X2=0 $Y2=0
cc_202 D N_A_215_367#_M1000_g 2.10277e-19 $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_203 N_D_c_273_n N_A_215_367#_c_320_n 0.006606f $X=2.505 $Y=0.955 $X2=0 $Y2=0
cc_204 N_D_M1011_g N_A_215_367#_c_320_n 0.00703575f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_D_c_273_n N_A_215_367#_c_321_n 0.00955838f $X=2.505 $Y=0.955 $X2=0
+ $Y2=0
cc_206 N_D_M1007_g N_A_215_367#_c_322_n 0.010995f $X=2.8 $Y=2.045 $X2=0 $Y2=0
cc_207 D N_A_215_367#_c_322_n 0.0186925f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_208 N_D_c_278_n N_A_215_367#_c_322_n 8.0758e-19 $X=2.8 $Y=2.79 $X2=0 $Y2=0
cc_209 N_D_c_273_n N_A_215_367#_c_323_n 0.00512959f $X=2.505 $Y=0.955 $X2=0
+ $Y2=0
cc_210 N_D_M1007_g N_A_215_367#_c_323_n 0.0116727f $X=2.8 $Y=2.045 $X2=0 $Y2=0
cc_211 N_D_c_273_n N_A_215_367#_c_324_n 0.0213197f $X=2.505 $Y=0.955 $X2=0 $Y2=0
cc_212 N_D_c_273_n N_A_215_367#_c_326_n 0.00547566f $X=2.505 $Y=0.955 $X2=0
+ $Y2=0
cc_213 N_D_M1007_g N_A_215_367#_c_326_n 0.00244062f $X=2.8 $Y=2.045 $X2=0 $Y2=0
cc_214 N_D_c_273_n N_A_215_367#_c_327_n 0.0054365f $X=2.505 $Y=0.955 $X2=0 $Y2=0
cc_215 N_D_M1011_g N_A_215_367#_c_327_n 0.00399102f $X=2.505 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_D_M1007_g N_VPWR_c_418_n 0.00165094f $X=2.8 $Y=2.045 $X2=0 $Y2=0
cc_217 D N_VPWR_c_418_n 0.0557897f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_218 N_D_c_278_n N_VPWR_c_418_n 0.00812811f $X=2.8 $Y=2.79 $X2=0 $Y2=0
cc_219 N_D_M1007_g N_VPWR_c_419_n 0.00817374f $X=2.8 $Y=2.045 $X2=0 $Y2=0
cc_220 D N_VPWR_c_419_n 0.0515111f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_221 D N_VPWR_c_423_n 0.010639f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_222 N_D_c_278_n N_VPWR_c_423_n 0.0052824f $X=2.8 $Y=2.79 $X2=0 $Y2=0
cc_223 D N_VPWR_c_416_n 0.0100383f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_224 N_D_c_278_n N_VPWR_c_416_n 0.00386935f $X=2.8 $Y=2.79 $X2=0 $Y2=0
cc_225 N_D_c_273_n N_VGND_c_483_n 6.13024e-19 $X=2.505 $Y=0.955 $X2=0 $Y2=0
cc_226 N_D_M1011_g N_VGND_c_483_n 0.00536427f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_227 N_D_c_273_n N_VGND_c_485_n 0.00517774f $X=2.505 $Y=0.955 $X2=0 $Y2=0
cc_228 N_D_M1011_g N_VGND_c_485_n 0.0183505f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_229 N_D_M1011_g N_VGND_c_487_n 0.00449212f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A_215_367#_c_331_n N_VPWR_c_418_n 0.0148223f $X=1.32 $Y=1.96 $X2=0
+ $Y2=0
cc_231 N_A_215_367#_M1000_g N_VPWR_c_419_n 0.0180379f $X=3.325 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_A_215_367#_M1000_g N_VPWR_c_420_n 0.00361735f $X=3.325 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_215_367#_c_322_n N_VPWR_c_420_n 0.0118805f $X=2.585 $Y=1.96 $X2=0
+ $Y2=0
cc_234 N_A_215_367#_c_323_n N_VPWR_c_420_n 0.0206321f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_235 N_A_215_367#_c_324_n N_VPWR_c_420_n 0.00361785f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_236 N_A_215_367#_M1000_g N_VPWR_c_424_n 0.00525069f $X=3.325 $Y=2.465 $X2=0
+ $Y2=0
cc_237 N_A_215_367#_M1000_g N_VPWR_c_416_n 0.00983341f $X=3.325 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A_215_367#_c_327_n X 0.00428002f $X=3.25 $Y=1.185 $X2=0 $Y2=0
cc_239 N_A_215_367#_M1000_g X 0.0115027f $X=3.325 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_215_367#_c_323_n X 0.0269573f $X=3.25 $Y=1.35 $X2=0 $Y2=0
cc_241 N_A_215_367#_c_324_n X 0.00824344f $X=3.25 $Y=1.35 $X2=0 $Y2=0
cc_242 N_A_215_367#_c_327_n X 0.006396f $X=3.25 $Y=1.185 $X2=0 $Y2=0
cc_243 N_A_215_367#_M1000_g X 0.00339266f $X=3.325 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A_215_367#_c_327_n N_X_c_464_n 0.0061838f $X=3.25 $Y=1.185 $X2=0 $Y2=0
cc_245 N_A_215_367#_c_317_n N_VGND_c_482_n 0.0181112f $X=1.375 $Y=0.485 $X2=0
+ $Y2=0
cc_246 N_A_215_367#_c_320_n N_VGND_c_483_n 0.0097297f $X=2.49 $Y=0.945 $X2=0
+ $Y2=0
cc_247 N_A_215_367#_c_323_n N_VGND_c_483_n 0.0215141f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_248 N_A_215_367#_c_324_n N_VGND_c_483_n 0.00238923f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_249 N_A_215_367#_c_317_n N_VGND_c_485_n 0.0280121f $X=1.375 $Y=0.485 $X2=0
+ $Y2=0
cc_250 N_A_215_367#_c_320_n N_VGND_c_485_n 0.00531576f $X=2.49 $Y=0.945 $X2=0
+ $Y2=0
cc_251 N_A_215_367#_c_323_n N_VGND_c_485_n 0.00658298f $X=3.25 $Y=1.35 $X2=0
+ $Y2=0
cc_252 N_A_215_367#_c_326_n N_VGND_c_485_n 0.00200959f $X=2.61 $Y=1.35 $X2=0
+ $Y2=0
cc_253 N_A_215_367#_c_327_n N_VGND_c_485_n 0.00434805f $X=3.25 $Y=1.185 $X2=0
+ $Y2=0
cc_254 N_A_215_367#_c_327_n N_VGND_c_486_n 0.0054895f $X=3.25 $Y=1.185 $X2=0
+ $Y2=0
cc_255 N_A_215_367#_M1001_s N_VGND_c_487_n 0.00215176f $X=1.085 $Y=0.235 $X2=0
+ $Y2=0
cc_256 N_A_215_367#_c_317_n N_VGND_c_487_n 0.0170321f $X=1.375 $Y=0.485 $X2=0
+ $Y2=0
cc_257 N_A_215_367#_c_320_n N_VGND_c_487_n 0.0330477f $X=2.49 $Y=0.945 $X2=0
+ $Y2=0
cc_258 N_A_215_367#_c_327_n N_VGND_c_487_n 0.0114319f $X=3.25 $Y=1.185 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_416_n N_X_M1000_d 0.00336915f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_c_420_n X 0.048041f $X=3.065 $Y=1.98 $X2=0 $Y2=0
cc_261 N_VPWR_c_424_n X 0.0217502f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_262 N_VPWR_c_416_n X 0.0123631f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_263 N_X_c_464_n N_VGND_c_486_n 0.0257063f $X=3.525 $Y=0.405 $X2=0 $Y2=0
cc_264 N_X_M1006_d N_VGND_c_487_n 0.00215158f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_265 N_X_c_464_n N_VGND_c_487_n 0.0150959f $X=3.525 $Y=0.405 $X2=0 $Y2=0
cc_266 N_VGND_c_487_n A_300_47# 0.00303238f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_267 N_VGND_c_487_n A_372_47# 0.00314438f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_268 N_VGND_c_487_n A_444_47# 0.00314438f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
