* File: sky130_fd_sc_lp__nand4b_4.pex.spice
* Created: Wed Sep  2 10:06:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4B_4%A_N 3 7 9 13 16
c34 13 0 7.10529e-20 $X=0.27 $Y=1.46
r35 15 16 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=0.475 $Y=1.46
+ $X2=0.825 $Y2=1.46
r36 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.475 $Y2=1.46
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.46 $X2=0.27 $Y2=1.46
r38 9 13 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.46
r39 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.825 $Y=1.625
+ $X2=0.825 $Y2=1.46
r40 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.825 $Y=1.625
+ $X2=0.825 $Y2=2.465
r41 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=1.46
r42 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%A_27_51# 1 2 9 13 17 21 25 29 33 37 41 43
+ 44 47 49 52 60 63 64 74
c118 74 0 7.10529e-20 $X=2.715 $Y=1.51
r119 71 72 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.205 $Y=1.51
+ $X2=2.285 $Y2=1.51
r120 70 71 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=1.855 $Y=1.51
+ $X2=2.205 $Y2=1.51
r121 69 70 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.695 $Y=1.51
+ $X2=1.855 $Y2=1.51
r122 68 69 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.425 $Y=1.51
+ $X2=1.695 $Y2=1.51
r123 61 74 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.635 $Y=1.51
+ $X2=2.715 $Y2=1.51
r124 61 72 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=2.635 $Y=1.51
+ $X2=2.285 $Y2=1.51
r125 60 61 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.635
+ $Y=1.51 $X2=2.635 $Y2=1.51
r126 58 68 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.275 $Y=1.51
+ $X2=1.425 $Y2=1.51
r127 58 65 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.275 $Y=1.51
+ $X2=1.265 $Y2=1.51
r128 57 60 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.275 $Y=1.51
+ $X2=2.635 $Y2=1.51
r129 57 58 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.275
+ $Y=1.51 $X2=1.275 $Y2=1.51
r130 55 64 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.855 $Y=1.51
+ $X2=0.73 $Y2=1.51
r131 55 57 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.855 $Y=1.51
+ $X2=1.275 $Y2=1.51
r132 53 64 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.69 $Y=1.595
+ $X2=0.73 $Y2=1.51
r133 53 63 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=1.595
+ $X2=0.69 $Y2=1.93
r134 52 64 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.425
+ $X2=0.73 $Y2=1.51
r135 51 52 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=0.73 $Y=1.195
+ $X2=0.73 $Y2=1.425
r136 47 63 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=2.095
+ $X2=0.61 $Y2=1.93
r137 47 49 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=0.61 $Y=2.095
+ $X2=0.61 $Y2=2.91
r138 43 51 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.605 $Y=1.11
+ $X2=0.73 $Y2=1.195
r139 43 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.11
+ $X2=0.345 $Y2=1.11
r140 39 44 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=1.025
+ $X2=0.345 $Y2=1.11
r141 39 41 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=0.22 $Y=1.025
+ $X2=0.22 $Y2=0.42
r142 35 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.345
+ $X2=2.715 $Y2=1.51
r143 35 37 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.715 $Y=1.345
+ $X2=2.715 $Y2=0.675
r144 31 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.675
+ $X2=2.635 $Y2=1.51
r145 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.635 $Y=1.675
+ $X2=2.635 $Y2=2.465
r146 27 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.345
+ $X2=2.285 $Y2=1.51
r147 27 29 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.285 $Y=1.345
+ $X2=2.285 $Y2=0.675
r148 23 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.675
+ $X2=2.205 $Y2=1.51
r149 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.205 $Y=1.675
+ $X2=2.205 $Y2=2.465
r150 19 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=1.51
r151 19 21 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=0.675
r152 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.675
+ $X2=1.695 $Y2=1.51
r153 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.695 $Y=1.675
+ $X2=1.695 $Y2=2.465
r154 11 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.51
r155 11 13 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=0.675
r156 7 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.675
+ $X2=1.265 $Y2=1.51
r157 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.265 $Y=1.675
+ $X2=1.265 $Y2=2.465
r158 2 49 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.485
+ $Y=1.835 $X2=0.61 $Y2=2.91
r159 2 47 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.485
+ $Y=1.835 $X2=0.61 $Y2=2.095
r160 1 41 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.255 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%B 3 7 11 15 19 23 27 31 38 39 59 62 68
r81 60 62 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=4.535 $Y=1.602
+ $X2=4.2 $Y2=1.602
r82 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=1.51 $X2=4.535 $Y2=1.51
r83 57 59 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.515 $Y=1.51
+ $X2=4.535 $Y2=1.51
r84 56 57 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.375 $Y=1.51
+ $X2=4.515 $Y2=1.51
r85 55 62 0.162316 $w=3.53e-07 $l=5e-09 $layer=LI1_cond $X=4.195 $Y=1.602
+ $X2=4.2 $Y2=1.602
r86 54 56 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.195 $Y=1.51
+ $X2=4.375 $Y2=1.51
r87 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.195
+ $Y=1.51 $X2=4.195 $Y2=1.51
r88 52 54 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.085 $Y=1.51
+ $X2=4.195 $Y2=1.51
r89 51 52 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.945 $Y=1.51
+ $X2=4.085 $Y2=1.51
r90 50 68 3.11953 $w=3.53e-07 $l=1e-08 $layer=LI1_cond $X=3.855 $Y=1.602
+ $X2=3.845 $Y2=1.602
r91 49 51 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=1.51
+ $X2=3.945 $Y2=1.51
r92 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.855
+ $Y=1.51 $X2=3.855 $Y2=1.51
r93 47 49 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=3.655 $Y=1.51
+ $X2=3.855 $Y2=1.51
r94 46 47 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.515 $Y=1.51
+ $X2=3.655 $Y2=1.51
r95 42 44 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.085 $Y=1.51
+ $X2=3.145 $Y2=1.51
r96 39 60 0.81158 $w=3.53e-07 $l=2.5e-08 $layer=LI1_cond $X=4.56 $Y=1.602
+ $X2=4.535 $Y2=1.602
r97 38 55 3.73327 $w=3.53e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.602
+ $X2=4.195 $Y2=1.602
r98 38 50 7.30422 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=4.08 $Y=1.602
+ $X2=3.855 $Y2=1.602
r99 36 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.175 $Y=1.51
+ $X2=3.515 $Y2=1.51
r100 36 44 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.175 $Y=1.51
+ $X2=3.145 $Y2=1.51
r101 35 68 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.175 $Y=1.515
+ $X2=3.845 $Y2=1.515
r102 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.175
+ $Y=1.51 $X2=3.175 $Y2=1.51
r103 29 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.515 $Y=1.345
+ $X2=4.515 $Y2=1.51
r104 29 31 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.515 $Y=1.345
+ $X2=4.515 $Y2=0.675
r105 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.675
+ $X2=4.375 $Y2=1.51
r106 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.375 $Y=1.675
+ $X2=4.375 $Y2=2.465
r107 21 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.085 $Y=1.345
+ $X2=4.085 $Y2=1.51
r108 21 23 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.085 $Y=1.345
+ $X2=4.085 $Y2=0.675
r109 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.675
+ $X2=3.945 $Y2=1.51
r110 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.945 $Y=1.675
+ $X2=3.945 $Y2=2.465
r111 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.345
+ $X2=3.655 $Y2=1.51
r112 13 15 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.655 $Y=1.345
+ $X2=3.655 $Y2=0.675
r113 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.675
+ $X2=3.515 $Y2=1.51
r114 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.515 $Y=1.675
+ $X2=3.515 $Y2=2.465
r115 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.345
+ $X2=3.145 $Y2=1.51
r116 5 7 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.145 $Y=1.345
+ $X2=3.145 $Y2=0.675
r117 1 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.675
+ $X2=3.085 $Y2=1.51
r118 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.085 $Y=1.675
+ $X2=3.085 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%C 3 7 11 15 19 23 27 31 33 34 58 59 61 73
r88 61 73 2.7304 $w=3.23e-07 $l=7.7e-08 $layer=LI1_cond $X=5.923 $Y=1.587 $X2=6
+ $Y2=1.587
r89 57 59 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.755 $Y=1.51
+ $X2=6.855 $Y2=1.51
r90 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.755
+ $Y=1.51 $X2=6.755 $Y2=1.51
r91 55 57 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=6.435 $Y=1.51
+ $X2=6.755 $Y2=1.51
r92 54 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.345 $Y=1.51
+ $X2=6.435 $Y2=1.51
r93 52 54 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.075 $Y=1.51
+ $X2=6.345 $Y2=1.51
r94 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.075
+ $Y=1.51 $X2=6.075 $Y2=1.51
r95 50 52 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.005 $Y=1.51
+ $X2=6.075 $Y2=1.51
r96 49 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.915 $Y=1.51
+ $X2=6.005 $Y2=1.51
r97 47 49 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.735 $Y=1.51
+ $X2=5.915 $Y2=1.51
r98 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.735
+ $Y=1.51 $X2=5.735 $Y2=1.51
r99 45 47 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.575 $Y=1.51
+ $X2=5.735 $Y2=1.51
r100 44 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.485 $Y=1.51
+ $X2=5.575 $Y2=1.51
r101 42 44 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.395 $Y=1.51
+ $X2=5.485 $Y2=1.51
r102 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.395
+ $Y=1.51 $X2=5.395 $Y2=1.51
r103 39 42 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.145 $Y=1.51
+ $X2=5.395 $Y2=1.51
r104 34 53 2.9639 $w=3.23e-07 $l=1e-08 $layer=LI1_cond $X=6.085 $Y=1.587
+ $X2=6.075 $Y2=1.587
r105 34 53 2.51764 $w=3.23e-07 $l=7.1e-08 $layer=LI1_cond $X=6.004 $Y=1.587
+ $X2=6.075 $Y2=1.587
r106 34 73 0.141839 $w=3.23e-07 $l=4e-09 $layer=LI1_cond $X=6.004 $Y=1.587 $X2=6
+ $Y2=1.587
r107 34 58 40.2596 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=6.085 $Y=1.51
+ $X2=6.755 $Y2=1.51
r108 34 61 0.141839 $w=3.23e-07 $l=4e-09 $layer=LI1_cond $X=5.919 $Y=1.587
+ $X2=5.923 $Y2=1.587
r109 34 48 6.5246 $w=3.23e-07 $l=1.84e-07 $layer=LI1_cond $X=5.919 $Y=1.587
+ $X2=5.735 $Y2=1.587
r110 33 48 7.62385 $w=3.23e-07 $l=2.15e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.735 $Y2=1.587
r111 33 43 4.43247 $w=3.23e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.395 $Y2=1.587
r112 29 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.855 $Y=1.345
+ $X2=6.855 $Y2=1.51
r113 29 31 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.855 $Y=1.345
+ $X2=6.855 $Y2=0.745
r114 25 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.435 $Y=1.675
+ $X2=6.435 $Y2=1.51
r115 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.435 $Y=1.675
+ $X2=6.435 $Y2=2.465
r116 21 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.345
+ $X2=6.345 $Y2=1.51
r117 21 23 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.345 $Y=1.345
+ $X2=6.345 $Y2=0.745
r118 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.005 $Y=1.675
+ $X2=6.005 $Y2=1.51
r119 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.005 $Y=1.675
+ $X2=6.005 $Y2=2.465
r120 13 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.345
+ $X2=5.915 $Y2=1.51
r121 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.915 $Y=1.345
+ $X2=5.915 $Y2=0.745
r122 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.675
+ $X2=5.575 $Y2=1.51
r123 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.575 $Y=1.675
+ $X2=5.575 $Y2=2.465
r124 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=1.345
+ $X2=5.485 $Y2=1.51
r125 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.485 $Y=1.345 $X2=5.485
+ $Y2=0.745
r126 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.675
+ $X2=5.145 $Y2=1.51
r127 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.145 $Y=1.675
+ $X2=5.145 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%D 3 7 11 15 19 23 27 31 38 39 40 57 61 70
c80 57 0 1.40803e-19 $X=8.575 $Y=1.51
c81 11 0 5.39005e-20 $X=7.665 $Y=2.465
c82 7 0 1.32946e-19 $X=7.285 $Y=0.745
c83 3 0 1.51739e-19 $X=7.235 $Y=2.465
r84 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.735
+ $Y=1.51 $X2=8.735 $Y2=1.51
r85 57 59 23.8025 $w=3.24e-07 $l=1.6e-07 $layer=POLY_cond $X=8.575 $Y=1.51
+ $X2=8.735 $Y2=1.51
r86 56 57 7.43827 $w=3.24e-07 $l=5e-08 $layer=POLY_cond $X=8.525 $Y=1.51
+ $X2=8.575 $Y2=1.51
r87 55 61 10.106 $w=3.23e-07 $l=2.85e-07 $layer=LI1_cond $X=8.395 $Y=1.587
+ $X2=8.11 $Y2=1.587
r88 54 56 19.3395 $w=3.24e-07 $l=1.3e-07 $layer=POLY_cond $X=8.395 $Y=1.51
+ $X2=8.525 $Y2=1.51
r89 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.395
+ $Y=1.51 $X2=8.395 $Y2=1.51
r90 52 54 37.1914 $w=3.24e-07 $l=2.5e-07 $layer=POLY_cond $X=8.145 $Y=1.51
+ $X2=8.395 $Y2=1.51
r91 51 52 7.43827 $w=3.24e-07 $l=5e-08 $layer=POLY_cond $X=8.095 $Y=1.51
+ $X2=8.145 $Y2=1.51
r92 50 61 1.95029 $w=3.23e-07 $l=5.5e-08 $layer=LI1_cond $X=8.055 $Y=1.587
+ $X2=8.11 $Y2=1.587
r93 49 51 5.95062 $w=3.24e-07 $l=4e-08 $layer=POLY_cond $X=8.055 $Y=1.51
+ $X2=8.095 $Y2=1.51
r94 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.055
+ $Y=1.51 $X2=8.055 $Y2=1.51
r95 45 46 56.5309 $w=3.24e-07 $l=3.8e-07 $layer=POLY_cond $X=7.285 $Y=1.51
+ $X2=7.665 $Y2=1.51
r96 44 45 7.43827 $w=3.24e-07 $l=5e-08 $layer=POLY_cond $X=7.235 $Y=1.51
+ $X2=7.285 $Y2=1.51
r97 40 60 5.14167 $w=3.23e-07 $l=1.45e-07 $layer=LI1_cond $X=8.88 $Y=1.587
+ $X2=8.735 $Y2=1.587
r98 39 60 11.879 $w=3.23e-07 $l=3.35e-07 $layer=LI1_cond $X=8.4 $Y=1.587
+ $X2=8.735 $Y2=1.587
r99 39 55 0.177299 $w=3.23e-07 $l=5e-09 $layer=LI1_cond $X=8.4 $Y=1.587
+ $X2=8.395 $Y2=1.587
r100 38 50 4.78707 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=1.587
+ $X2=8.055 $Y2=1.587
r101 38 70 7.39638 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=1.587
+ $X2=7.785 $Y2=1.587
r102 36 49 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=7.715 $Y=1.51
+ $X2=8.055 $Y2=1.51
r103 36 46 7.43827 $w=3.24e-07 $l=5e-08 $layer=POLY_cond $X=7.715 $Y=1.51
+ $X2=7.665 $Y2=1.51
r104 35 70 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.715 $Y=1.51
+ $X2=7.785 $Y2=1.51
r105 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.715
+ $Y=1.51 $X2=7.715 $Y2=1.51
r106 29 57 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.575 $Y=1.345
+ $X2=8.575 $Y2=1.51
r107 29 31 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.575 $Y=1.345
+ $X2=8.575 $Y2=0.745
r108 25 56 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.525 $Y=1.675
+ $X2=8.525 $Y2=1.51
r109 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.525 $Y=1.675
+ $X2=8.525 $Y2=2.465
r110 21 52 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.145 $Y=1.345
+ $X2=8.145 $Y2=1.51
r111 21 23 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.145 $Y=1.345
+ $X2=8.145 $Y2=0.745
r112 17 51 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=1.675
+ $X2=8.095 $Y2=1.51
r113 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.095 $Y=1.675
+ $X2=8.095 $Y2=2.465
r114 13 36 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.715 $Y=1.345
+ $X2=7.715 $Y2=1.51
r115 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.715 $Y=1.345
+ $X2=7.715 $Y2=0.745
r116 9 46 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=1.675
+ $X2=7.665 $Y2=1.51
r117 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.665 $Y=1.675
+ $X2=7.665 $Y2=2.465
r118 5 45 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.285 $Y=1.345
+ $X2=7.285 $Y2=1.51
r119 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.285 $Y=1.345 $X2=7.285
+ $Y2=0.745
r120 1 44 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.235 $Y=1.675
+ $X2=7.235 $Y2=1.51
r121 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.235 $Y=1.675
+ $X2=7.235 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%VPWR 1 2 3 4 5 6 7 8 9 30 36 42 46 50 54 58
+ 62 68 70 72 77 78 80 81 82 83 85 86 87 99 108 112 117 123 126 129 132 136
r146 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r147 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r150 121 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r151 121 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r152 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r153 118 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=7.88 $Y2=3.33
r154 118 120 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 117 135 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.847 $Y2=3.33
r156 117 120 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.4 $Y2=3.33
r157 116 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r158 116 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r159 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r160 113 129 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=7.185 $Y=3.33
+ $X2=6.89 $Y2=3.33
r161 113 115 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.185 $Y=3.33
+ $X2=7.44 $Y2=3.33
r162 112 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.88 $Y2=3.33
r163 112 115 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r164 111 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r165 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r166 108 129 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.89 $Y2=3.33
r167 108 110 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 107 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r169 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r170 104 126 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=4.76 $Y2=3.33
r171 104 106 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=5.52 $Y2=3.33
r172 103 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r173 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r174 100 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=3.73 $Y2=3.33
r175 100 102 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=4.08 $Y2=3.33
r176 99 126 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.76 $Y2=3.33
r177 99 102 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r178 98 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r179 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r180 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r181 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r182 91 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r183 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 87 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r185 87 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r186 87 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r187 85 106 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.625 $Y=3.33
+ $X2=5.52 $Y2=3.33
r188 85 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.625 $Y=3.33
+ $X2=5.79 $Y2=3.33
r189 84 110 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.955 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 84 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.955 $Y=3.33
+ $X2=5.79 $Y2=3.33
r191 82 97 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 82 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.85 $Y2=3.33
r193 80 94 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.68 $Y2=3.33
r194 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.95 $Y2=3.33
r195 79 97 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.64 $Y2=3.33
r196 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.95 $Y2=3.33
r197 77 90 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.72 $Y2=3.33
r198 77 78 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.06 $Y2=3.33
r199 76 94 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.68 $Y2=3.33
r200 76 78 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.06 $Y2=3.33
r201 72 75 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=8.74 $Y=2.005
+ $X2=8.74 $Y2=2.95
r202 70 135 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=8.74 $Y=3.245
+ $X2=8.847 $Y2=3.33
r203 70 75 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.74 $Y=3.245
+ $X2=8.74 $Y2=2.95
r204 66 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=3.33
r205 66 68 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=2.355
r206 62 65 14.1908 $w=5.88e-07 $l=7e-07 $layer=LI1_cond $X=6.89 $Y=2.27 $X2=6.89
+ $Y2=2.97
r207 60 129 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=3.245
+ $X2=6.89 $Y2=3.33
r208 60 65 5.57494 $w=5.88e-07 $l=2.75e-07 $layer=LI1_cond $X=6.89 $Y=3.245
+ $X2=6.89 $Y2=2.97
r209 56 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.79 $Y=3.245
+ $X2=5.79 $Y2=3.33
r210 56 58 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=5.79 $Y=3.245
+ $X2=5.79 $Y2=2.375
r211 52 126 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=3.245
+ $X2=4.76 $Y2=3.33
r212 52 54 15.5312 $w=6.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.76 $Y=3.245
+ $X2=4.76 $Y2=2.375
r213 48 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=3.245
+ $X2=3.73 $Y2=3.33
r214 48 50 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.73 $Y=3.245
+ $X2=3.73 $Y2=2.375
r215 47 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=3.33
+ $X2=2.85 $Y2=3.33
r216 46 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=3.33
+ $X2=3.73 $Y2=3.33
r217 46 47 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.565 $Y=3.33
+ $X2=3.015 $Y2=3.33
r218 42 45 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.85 $Y=2.2
+ $X2=2.85 $Y2=2.97
r219 40 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=3.33
r220 40 45 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=2.97
r221 36 39 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.95 $Y=2.21
+ $X2=1.95 $Y2=2.97
r222 34 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=3.33
r223 34 39 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=2.97
r224 30 33 48.603 $w=2.28e-07 $l=9.7e-07 $layer=LI1_cond $X=1.06 $Y=1.98
+ $X2=1.06 $Y2=2.95
r225 28 78 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=3.33
r226 28 33 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=2.95
r227 9 75 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.6
+ $Y=1.835 $X2=8.74 $Y2=2.95
r228 9 72 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=8.6
+ $Y=1.835 $X2=8.74 $Y2=2.005
r229 8 68 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=7.74
+ $Y=1.835 $X2=7.88 $Y2=2.355
r230 7 65 200 $w=1.7e-07 $l=1.21704e-06 $layer=licon1_PDIFF $count=3 $X=6.51
+ $Y=1.835 $X2=6.68 $Y2=2.97
r231 7 62 200 $w=1.7e-07 $l=5.13006e-07 $layer=licon1_PDIFF $count=3 $X=6.51
+ $Y=1.835 $X2=6.68 $Y2=2.27
r232 6 58 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=5.65
+ $Y=1.835 $X2=5.79 $Y2=2.375
r233 5 54 150 $w=1.7e-07 $l=7.42159e-07 $layer=licon1_PDIFF $count=4 $X=4.45
+ $Y=1.835 $X2=4.93 $Y2=2.375
r234 4 50 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=3.59
+ $Y=1.835 $X2=3.73 $Y2=2.375
r235 3 45 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=2.97
r236 3 42 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=2.2
r237 2 39 400 $w=1.7e-07 $l=1.22169e-06 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.835 $X2=1.95 $Y2=2.97
r238 2 36 400 $w=1.7e-07 $l=4.56207e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.835 $X2=1.95 $Y2=2.21
r239 1 33 400 $w=1.7e-07 $l=1.18763e-06 $layer=licon1_PDIFF $count=1 $X=0.9
+ $Y=1.835 $X2=1.05 $Y2=2.95
r240 1 30 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.9
+ $Y=1.835 $X2=1.05 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%Y 1 2 3 4 5 6 7 8 9 10 33 39 41 42 43 44 47
+ 53 57 61 64 65 67 69 73 75 77 79 81 82 85 88 91 94 102 103 104 105 106 117 119
+ 123 128 134 139
c166 94 0 1.51739e-19 $X=7.485 $Y=1.85
c167 69 0 5.39005e-20 $X=7.355 $Y=1.85
r168 126 128 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=5.455 $Y=2.02
+ $X2=5.52 $Y2=2.02
r169 105 123 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.36 $Y=2.02
+ $X2=5.265 $Y2=2.02
r170 105 126 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.36 $Y=2.02
+ $X2=5.455 $Y2=2.02
r171 105 139 41.8466 $w=2.08e-07 $l=7.9e-07 $layer=LI1_cond $X=5.36 $Y=2.12
+ $X2=5.36 $Y2=2.91
r172 105 106 26.0636 $w=1.98e-07 $l=4.7e-07 $layer=LI1_cond $X=5.53 $Y=2.02
+ $X2=6 $Y2=2.02
r173 105 128 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=5.53 $Y=2.02
+ $X2=5.52 $Y2=2.02
r174 104 119 4.81226 $w=1.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=4.965 $Y=2.02
+ $X2=4.88 $Y2=2.035
r175 104 124 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=2.02
+ $X2=5.05 $Y2=2.02
r176 104 123 9.87091 $w=1.98e-07 $l=1.78e-07 $layer=LI1_cond $X=5.087 $Y=2.02
+ $X2=5.265 $Y2=2.02
r177 104 124 2.05182 $w=1.98e-07 $l=3.7e-08 $layer=LI1_cond $X=5.087 $Y=2.02
+ $X2=5.05 $Y2=2.02
r178 103 119 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.56 $Y=2.035
+ $X2=4.88 $Y2=2.035
r179 103 120 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.56 $Y=2.035
+ $X2=4.255 $Y2=2.035
r180 102 117 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.16 $Y=2.035
+ $X2=4.065 $Y2=2.035
r181 102 120 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.16 $Y=2.035
+ $X2=4.255 $Y2=2.035
r182 102 134 32.764 $w=2.88e-07 $l=7.9e-07 $layer=LI1_cond $X=4.16 $Y=2.12
+ $X2=4.16 $Y2=2.91
r183 102 117 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.03 $Y=2.035
+ $X2=4.065 $Y2=2.035
r184 98 99 4.86943 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=2.015
+ $X2=7.485 $Y2=2.1
r185 97 98 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=7.485 $Y=1.98
+ $X2=7.485 $Y2=2.015
r186 94 97 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=7.485 $Y=1.85
+ $X2=7.485 $Y2=1.98
r187 91 106 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=6.125 $Y=2.02
+ $X2=6 $Y2=2.02
r188 90 93 0.753086 $w=2.43e-07 $l=1.5e-08 $layer=LI1_cond $X=6.275 $Y=2.02
+ $X2=6.275 $Y2=2.035
r189 90 91 1.87978 $w=2e-07 $l=1.5e-07 $layer=LI1_cond $X=6.275 $Y=2.02
+ $X2=6.125 $Y2=2.02
r190 89 90 8.53498 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=6.275 $Y=1.85
+ $X2=6.275 $Y2=2.02
r191 88 102 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=4.03 $Y2=2.035
r192 87 88 15.3273 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.3 $Y=1.947
+ $X2=3.67 $Y2=1.947
r193 84 87 0.334041 $w=3.43e-07 $l=1e-08 $layer=LI1_cond $X=3.29 $Y=1.947
+ $X2=3.3 $Y2=1.947
r194 84 85 6.47515 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=3.29 $Y=1.947
+ $X2=3.185 $Y2=1.947
r195 77 101 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.31 $Y=2.1
+ $X2=8.31 $Y2=2.015
r196 77 79 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=8.31 $Y=2.1
+ $X2=8.31 $Y2=2.91
r197 76 98 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.615 $Y=2.015
+ $X2=7.485 $Y2=2.015
r198 75 101 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.215 $Y=2.015
+ $X2=8.31 $Y2=2.015
r199 75 76 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.215 $Y=2.015
+ $X2=7.615 $Y2=2.015
r200 73 99 21.5657 $w=1.78e-07 $l=3.5e-07 $layer=LI1_cond $X=7.445 $Y=2.45
+ $X2=7.445 $Y2=2.1
r201 70 89 2.8297 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.425 $Y=1.85
+ $X2=6.275 $Y2=1.85
r202 69 94 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.355 $Y=1.85
+ $X2=7.485 $Y2=1.85
r203 69 70 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=7.355 $Y=1.85
+ $X2=6.425 $Y2=1.85
r204 65 93 3.93284 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.275 $Y=2.12
+ $X2=6.275 $Y2=2.035
r205 65 67 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=6.275 $Y=2.12
+ $X2=6.275 $Y2=2.475
r206 64 104 1.64875 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.965 $Y=1.92
+ $X2=4.965 $Y2=2.02
r207 63 64 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.965 $Y=1.255
+ $X2=4.965 $Y2=1.92
r208 59 84 3.64154 $w=2.1e-07 $l=1.73e-07 $layer=LI1_cond $X=3.29 $Y=2.12
+ $X2=3.29 $Y2=1.947
r209 59 61 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=3.29 $Y=2.12
+ $X2=3.29 $Y2=2.46
r210 58 82 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.595 $Y=1.165
+ $X2=2.5 $Y2=1.165
r211 57 63 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.88 $Y=1.165
+ $X2=4.965 $Y2=1.255
r212 57 58 140.793 $w=1.78e-07 $l=2.285e-06 $layer=LI1_cond $X=4.88 $Y=1.165
+ $X2=2.595 $Y2=1.165
r213 56 81 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.515 $Y=1.86
+ $X2=2.4 $Y2=1.86
r214 56 85 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.515 $Y=1.86
+ $X2=3.185 $Y2=1.86
r215 51 82 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.5 $Y=1.075 $X2=2.5
+ $Y2=1.165
r216 51 53 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.5 $Y=1.075
+ $X2=2.5 $Y2=0.76
r217 47 49 46.5988 $w=2.28e-07 $l=9.3e-07 $layer=LI1_cond $X=2.4 $Y=1.98 $X2=2.4
+ $Y2=2.91
r218 45 81 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=1.945
+ $X2=2.4 $Y2=1.86
r219 45 47 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.4 $Y=1.945
+ $X2=2.4 $Y2=1.98
r220 43 82 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.405 $Y=1.165
+ $X2=2.5 $Y2=1.165
r221 43 44 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.405 $Y=1.165
+ $X2=1.735 $Y2=1.165
r222 41 81 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.285 $Y=1.86
+ $X2=2.4 $Y2=1.86
r223 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.285 $Y=1.86
+ $X2=1.615 $Y2=1.86
r224 37 44 6.92652 $w=1.8e-07 $l=1.51456e-07 $layer=LI1_cond $X=1.622 $Y=1.075
+ $X2=1.735 $Y2=1.165
r225 37 39 16.1342 $w=2.23e-07 $l=3.15e-07 $layer=LI1_cond $X=1.622 $Y=1.075
+ $X2=1.622 $Y2=0.76
r226 33 35 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.48 $Y=1.98
+ $X2=1.48 $Y2=2.91
r227 31 42 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.48 $Y=1.945
+ $X2=1.615 $Y2=1.86
r228 31 33 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.48 $Y=1.945
+ $X2=1.48 $Y2=1.98
r229 10 101 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=8.17
+ $Y=1.835 $X2=8.31 $Y2=2.095
r230 10 79 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.17
+ $Y=1.835 $X2=8.31 $Y2=2.91
r231 9 97 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=1.835 $X2=7.45 $Y2=1.98
r232 9 73 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=7.31
+ $Y=1.835 $X2=7.45 $Y2=2.45
r233 8 93 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=6.08
+ $Y=1.835 $X2=6.22 $Y2=2.035
r234 8 67 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=6.08
+ $Y=1.835 $X2=6.22 $Y2=2.475
r235 7 105 400 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.835 $X2=5.36 $Y2=2.115
r236 7 139 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.835 $X2=5.36 $Y2=2.91
r237 6 102 400 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=2.115
r238 6 134 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.16 $Y2=2.91
r239 5 87 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=1.835 $X2=3.3 $Y2=1.98
r240 5 61 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=3.16
+ $Y=1.835 $X2=3.3 $Y2=2.46
r241 4 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=2.91
r242 4 47 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=1.98
r243 3 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=1.835 $X2=1.48 $Y2=2.91
r244 3 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=1.835 $X2=1.48 $Y2=1.98
r245 2 53 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.255 $X2=2.5 $Y2=0.76
r246 1 39 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.255 $X2=1.64 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48 51
+ 54
r92 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r93 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r94 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r96 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r97 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.525 $Y=0 $X2=8.36
+ $Y2=0
r98 42 44 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.525 $Y=0 $X2=8.88
+ $Y2=0
r99 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r100 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r101 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r102 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.5
+ $Y2=0
r103 38 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.92 $Y2=0
r104 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=0 $X2=8.36
+ $Y2=0
r105 37 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.195 $Y=0
+ $X2=7.92 $Y2=0
r106 36 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r107 35 36 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r108 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 32 35 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=6.96
+ $Y2=0
r110 32 33 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r111 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r112 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r113 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.5
+ $Y2=0
r114 29 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=6.96 $Y2=0
r115 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r116 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r117 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r118 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r119 22 36 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6.96
+ $Y2=0
r120 22 33 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r121 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=0.085
+ $X2=8.36 $Y2=0
r122 18 20 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=8.36 $Y=0.085
+ $X2=8.36 $Y2=0.45
r123 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.085 $X2=7.5
+ $Y2=0
r124 14 16 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0.45
r125 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r126 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.4
r127 3 20 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.325 $X2=8.36 $Y2=0.45
r128 2 16 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.36
+ $Y=0.325 $X2=7.5 $Y2=0.45
r129 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.255 $X2=0.69 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%A_217_51# 1 2 3 4 5 18 22 30 33 35 37
r61 28 30 38.1193 $w=2.58e-07 $l=8.6e-07 $layer=LI1_cond $X=3.87 $Y=0.385
+ $X2=4.73 $Y2=0.385
r62 26 37 7.25953 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=0.385
+ $X2=2.93 $Y2=0.385
r63 26 28 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=3.095 $Y=0.385
+ $X2=3.87 $Y2=0.385
r64 23 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0.34
+ $X2=2.07 $Y2=0.34
r65 22 37 7.25953 $w=2.15e-07 $l=1.86145e-07 $layer=LI1_cond $X=2.765 $Y=0.34
+ $X2=2.93 $Y2=0.385
r66 22 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.765 $Y=0.34
+ $X2=2.235 $Y2=0.34
r67 19 33 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.34 $Y=0.34
+ $X2=1.192 $Y2=0.34
r68 18 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0.34
+ $X2=2.07 $Y2=0.34
r69 18 19 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.905 $Y=0.34
+ $X2=1.34 $Y2=0.34
r70 5 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.59
+ $Y=0.255 $X2=4.73 $Y2=0.4
r71 4 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.255 $X2=3.87 $Y2=0.4
r72 3 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.79
+ $Y=0.255 $X2=2.93 $Y2=0.4
r73 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.255 $X2=2.07 $Y2=0.4
r74 1 33 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.255 $X2=1.21 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%A_644_51# 1 2 3 4 13 19 21 22 23 24 27 29
c46 23 0 1.32946e-19 $X=6.475 $Y=1.165
r47 25 27 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.64 $Y=1.075
+ $X2=6.64 $Y2=0.69
r48 23 25 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=6.475 $Y=1.165
+ $X2=6.64 $Y2=1.075
r49 23 24 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.475 $Y=1.165
+ $X2=5.795 $Y2=1.165
r50 22 24 7.14503 $w=1.8e-07 $l=1.72218e-07 $layer=LI1_cond $X=5.662 $Y=1.075
+ $X2=5.795 $Y2=1.165
r51 21 31 2.89663 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=5.662 $Y=0.905
+ $X2=5.662 $Y2=0.815
r52 21 22 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=5.662 $Y=0.905
+ $X2=5.662 $Y2=1.075
r53 19 31 4.2484 $w=1.8e-07 $l=1.32e-07 $layer=LI1_cond $X=5.53 $Y=0.815
+ $X2=5.662 $Y2=0.815
r54 19 29 65.6212 $w=1.78e-07 $l=1.065e-06 $layer=LI1_cond $X=5.53 $Y=0.815
+ $X2=4.465 $Y2=0.815
r55 15 18 45.05 $w=2.18e-07 $l=8.6e-07 $layer=LI1_cond $X=3.44 $Y=0.795 $X2=4.3
+ $Y2=0.795
r56 13 29 6.17723 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=4.355 $Y=0.795
+ $X2=4.465 $Y2=0.795
r57 13 18 2.88111 $w=2.18e-07 $l=5.5e-08 $layer=LI1_cond $X=4.355 $Y=0.795
+ $X2=4.3 $Y2=0.795
r58 4 27 91 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_NDIFF $count=2 $X=6.42
+ $Y=0.325 $X2=6.64 $Y2=0.69
r59 3 31 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.325 $X2=5.7 $Y2=0.89
r60 2 18 182 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_NDIFF $count=1 $X=4.16
+ $Y=0.255 $X2=4.3 $Y2=0.79
r61 1 15 182 $w=1.7e-07 $l=6.35551e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.255 $X2=3.44 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_4%A_1025_65# 1 2 3 4 5 16 22 28 29 32 34 38
+ 41 42
c65 29 0 1.40803e-19 $X=7.165 $Y=1.16
r66 36 38 26.8165 $w=2.58e-07 $l=6.05e-07 $layer=LI1_cond $X=8.825 $Y=1.075
+ $X2=8.825 $Y2=0.47
r67 35 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.025 $Y=1.16
+ $X2=7.93 $Y2=1.16
r68 34 36 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=8.695 $Y=1.16
+ $X2=8.825 $Y2=1.075
r69 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.695 $Y=1.16
+ $X2=8.025 $Y2=1.16
r70 30 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=1.075
+ $X2=7.93 $Y2=1.16
r71 30 32 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=7.93 $Y=1.075
+ $X2=7.93 $Y2=0.47
r72 28 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.835 $Y=1.16
+ $X2=7.93 $Y2=1.16
r73 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.835 $Y=1.16
+ $X2=7.165 $Y2=1.16
r74 25 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.07 $Y=1.075
+ $X2=7.165 $Y2=1.16
r75 25 27 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=7.07 $Y=1.075
+ $X2=7.07 $Y2=0.47
r76 24 27 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=7.07 $Y=0.435
+ $X2=7.07 $Y2=0.47
r77 23 41 6.67463 $w=2.4e-07 $l=1.92678e-07 $layer=LI1_cond $X=6.295 $Y=0.345
+ $X2=6.13 $Y2=0.405
r78 22 24 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=6.975 $Y=0.345
+ $X2=7.07 $Y2=0.435
r79 22 23 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.975 $Y=0.345
+ $X2=6.295 $Y2=0.345
r80 16 41 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=0.405
+ $X2=6.13 $Y2=0.405
r81 16 18 26.6983 $w=2.98e-07 $l=6.95e-07 $layer=LI1_cond $X=5.965 $Y=0.405
+ $X2=5.27 $Y2=0.405
r82 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.65
+ $Y=0.325 $X2=8.79 $Y2=0.47
r83 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.325 $X2=7.93 $Y2=0.47
r84 3 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.93
+ $Y=0.325 $X2=7.07 $Y2=0.47
r85 2 41 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.99
+ $Y=0.325 $X2=6.13 $Y2=0.45
r86 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.325 $X2=5.27 $Y2=0.45
.ends

