* File: sky130_fd_sc_lp__xnor2_lp.spice
* Created: Wed Sep  2 10:40:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor2_lp.pex.spice"
.subckt sky130_fd_sc_lp__xnor2_lp  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 N_A_112_92#_M1009_d N_A_82_66#_M1009_g N_Y_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.1155 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_112_92#_M1001_d N_B_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1155 PD=0.86 PS=1.39 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_112_92#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_510_125# N_A_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_82_66#_M1008_d N_B_M1008_g A_510_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_82_66#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1006 A_280_419# N_B_M1006_g N_Y_M1000_d VPB PHIGHVT L=0.25 W=1 AD=0.12 AS=0.14
+ PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_280_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1007 N_A_82_66#_M1007_d N_A_M1007_g N_VPWR_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_82_66#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.275 AS=0.14 PD=2.55 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__xnor2_lp.pxi.spice"
*
.ends
*
*
