* File: sky130_fd_sc_lp__dfxtp_2.pxi.spice
* Created: Wed Sep  2 09:45:14 2020
* 
x_PM_SKY130_FD_SC_LP__DFXTP_2%CLK N_CLK_c_158_n N_CLK_M1023_g N_CLK_M1021_g
+ N_CLK_c_160_n CLK CLK CLK CLK CLK N_CLK_c_162_n N_CLK_c_163_n
+ PM_SKY130_FD_SC_LP__DFXTP_2%CLK
x_PM_SKY130_FD_SC_LP__DFXTP_2%D N_D_M1012_g N_D_M1010_g D D N_D_c_183_n
+ N_D_c_184_n PM_SKY130_FD_SC_LP__DFXTP_2%D
x_PM_SKY130_FD_SC_LP__DFXTP_2%A_240_443# N_A_240_443#_M1009_s
+ N_A_240_443#_M1013_s N_A_240_443#_M1022_g N_A_240_443#_M1004_g
+ N_A_240_443#_M1018_g N_A_240_443#_c_225_n N_A_240_443#_c_235_n
+ N_A_240_443#_M1017_g N_A_240_443#_c_226_n N_A_240_443#_c_236_n
+ N_A_240_443#_c_227_n N_A_240_443#_c_238_n N_A_240_443#_c_239_n
+ N_A_240_443#_c_240_n N_A_240_443#_c_241_n N_A_240_443#_c_242_n
+ N_A_240_443#_c_228_n N_A_240_443#_c_229_n N_A_240_443#_c_245_n
+ N_A_240_443#_c_246_n N_A_240_443#_c_265_p N_A_240_443#_c_272_p
+ N_A_240_443#_c_230_n N_A_240_443#_c_231_n N_A_240_443#_c_248_n
+ N_A_240_443#_c_249_n N_A_240_443#_c_232_n
+ PM_SKY130_FD_SC_LP__DFXTP_2%A_240_443#
x_PM_SKY130_FD_SC_LP__DFXTP_2%A_679_93# N_A_679_93#_M1000_d N_A_679_93#_M1011_d
+ N_A_679_93#_M1024_g N_A_679_93#_M1005_g N_A_679_93#_c_386_n
+ N_A_679_93#_c_391_n N_A_679_93#_c_392_n N_A_679_93#_c_403_n
+ N_A_679_93#_c_387_n N_A_679_93#_c_388_n PM_SKY130_FD_SC_LP__DFXTP_2%A_679_93#
x_PM_SKY130_FD_SC_LP__DFXTP_2%A_551_119# N_A_551_119#_M1015_d
+ N_A_551_119#_M1022_d N_A_551_119#_M1011_g N_A_551_119#_M1000_g
+ N_A_551_119#_c_449_n N_A_551_119#_c_450_n N_A_551_119#_c_451_n
+ N_A_551_119#_c_452_n N_A_551_119#_c_453_n N_A_551_119#_c_454_n
+ PM_SKY130_FD_SC_LP__DFXTP_2%A_551_119#
x_PM_SKY130_FD_SC_LP__DFXTP_2%A_110_62# N_A_110_62#_M1023_d N_A_110_62#_M1021_d
+ N_A_110_62#_c_514_n N_A_110_62#_c_515_n N_A_110_62#_M1013_g
+ N_A_110_62#_M1009_g N_A_110_62#_c_528_n N_A_110_62#_c_529_n
+ N_A_110_62#_c_518_n N_A_110_62#_c_519_n N_A_110_62#_M1015_g
+ N_A_110_62#_c_521_n N_A_110_62#_M1002_g N_A_110_62#_c_531_n
+ N_A_110_62#_M1014_g N_A_110_62#_M1006_g N_A_110_62#_c_523_n
+ N_A_110_62#_c_524_n N_A_110_62#_c_533_n N_A_110_62#_c_525_n
+ N_A_110_62#_c_526_n PM_SKY130_FD_SC_LP__DFXTP_2%A_110_62#
x_PM_SKY130_FD_SC_LP__DFXTP_2%A_1175_93# N_A_1175_93#_M1003_d
+ N_A_1175_93#_M1007_d N_A_1175_93#_M1001_g N_A_1175_93#_c_644_n
+ N_A_1175_93#_M1020_g N_A_1175_93#_c_645_n N_A_1175_93#_M1016_g
+ N_A_1175_93#_M1008_g N_A_1175_93#_c_646_n N_A_1175_93#_c_647_n
+ N_A_1175_93#_M1025_g N_A_1175_93#_M1019_g N_A_1175_93#_c_649_n
+ N_A_1175_93#_c_650_n N_A_1175_93#_c_651_n N_A_1175_93#_c_652_n
+ N_A_1175_93#_c_663_n N_A_1175_93#_c_653_n N_A_1175_93#_c_664_n
+ N_A_1175_93#_c_654_n N_A_1175_93#_c_655_n
+ PM_SKY130_FD_SC_LP__DFXTP_2%A_1175_93#
x_PM_SKY130_FD_SC_LP__DFXTP_2%A_1004_379# N_A_1004_379#_M1018_d
+ N_A_1004_379#_M1014_d N_A_1004_379#_M1003_g N_A_1004_379#_M1007_g
+ N_A_1004_379#_c_747_n N_A_1004_379#_c_748_n N_A_1004_379#_c_740_n
+ N_A_1004_379#_c_741_n N_A_1004_379#_c_742_n N_A_1004_379#_c_743_n
+ N_A_1004_379#_c_744_n N_A_1004_379#_c_745_n
+ PM_SKY130_FD_SC_LP__DFXTP_2%A_1004_379#
x_PM_SKY130_FD_SC_LP__DFXTP_2%VPWR N_VPWR_M1021_s N_VPWR_M1013_d N_VPWR_M1005_d
+ N_VPWR_M1020_d N_VPWR_M1008_s N_VPWR_M1019_s N_VPWR_c_815_n N_VPWR_c_816_n
+ N_VPWR_c_817_n N_VPWR_c_818_n N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_821_n
+ N_VPWR_c_822_n N_VPWR_c_823_n N_VPWR_c_824_n VPWR N_VPWR_c_825_n
+ N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n N_VPWR_c_829_n N_VPWR_c_830_n
+ N_VPWR_c_831_n N_VPWR_c_814_n PM_SKY130_FD_SC_LP__DFXTP_2%VPWR
x_PM_SKY130_FD_SC_LP__DFXTP_2%A_432_119# N_A_432_119#_M1012_d
+ N_A_432_119#_M1010_d N_A_432_119#_c_914_n N_A_432_119#_c_915_n
+ N_A_432_119#_c_919_n N_A_432_119#_c_916_n
+ PM_SKY130_FD_SC_LP__DFXTP_2%A_432_119#
x_PM_SKY130_FD_SC_LP__DFXTP_2%Q N_Q_M1016_d N_Q_M1008_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DFXTP_2%Q
x_PM_SKY130_FD_SC_LP__DFXTP_2%VGND N_VGND_M1023_s N_VGND_M1009_d N_VGND_M1024_d
+ N_VGND_M1001_d N_VGND_M1016_s N_VGND_M1025_s N_VGND_c_961_n N_VGND_c_962_n
+ N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n
+ N_VGND_c_968_n N_VGND_c_969_n VGND N_VGND_c_970_n N_VGND_c_971_n
+ N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n N_VGND_c_975_n N_VGND_c_976_n
+ PM_SKY130_FD_SC_LP__DFXTP_2%VGND
cc_1 VNB N_CLK_c_158_n 0.0252782f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.313
cc_2 VNB N_CLK_M1021_g 0.00891274f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.72
cc_3 VNB N_CLK_c_160_n 0.0243916f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.51
cc_4 VNB CLK 0.0333978f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_CLK_c_162_n 0.025499f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.005
cc_6 VNB N_CLK_c_163_n 0.0251373f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.84
cc_7 VNB N_D_c_183_n 0.0577599f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_D_c_184_n 0.0161668f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_9 VNB N_A_240_443#_M1004_g 0.0282456f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A_240_443#_M1018_g 0.0237089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_240_443#_c_225_n 0.0115358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_240_443#_c_226_n 0.0293224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_240_443#_c_227_n 0.00898128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_240_443#_c_228_n 0.00210547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_240_443#_c_229_n 0.00960891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_240_443#_c_230_n 0.00429714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_240_443#_c_231_n 0.0014079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_240_443#_c_232_n 0.0542647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_679_93#_M1024_g 0.033894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_679_93#_c_386_n 0.00314312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_679_93#_c_387_n 0.0101786f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.84
cc_22 VNB N_A_679_93#_c_388_n 0.0345016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_551_119#_c_449_n 0.00402001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_551_119#_c_450_n 0.0201819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_551_119#_c_451_n 0.00334676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_551_119#_c_452_n 0.00165495f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.005
cc_27 VNB N_A_551_119#_c_453_n 0.0340539f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.005
cc_28 VNB N_A_551_119#_c_454_n 0.0183868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_110_62#_c_514_n 0.0223132f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.72
cc_30 VNB N_A_110_62#_c_515_n 0.0185408f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.72
cc_31 VNB N_A_110_62#_M1013_g 0.0143476f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_32 VNB N_A_110_62#_M1009_g 0.0367626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_110_62#_c_518_n 0.0602509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_110_62#_c_519_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_110_62#_M1015_g 0.038621f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.005
cc_36 VNB N_A_110_62#_c_521_n 0.214531f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_37 VNB N_A_110_62#_M1006_g 0.0350856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_110_62#_c_523_n 0.0140036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_110_62#_c_524_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_110_62#_c_525_n 0.0253727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_110_62#_c_526_n 0.0181401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1175_93#_M1001_g 0.0252773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1175_93#_c_644_n 0.0522052f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_44 VNB N_A_1175_93#_c_645_n 0.017504f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_45 VNB N_A_1175_93#_c_646_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.005
cc_46 VNB N_A_1175_93#_c_647_n 0.0192431f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.84
cc_47 VNB N_A_1175_93#_M1019_g 0.0127435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1175_93#_c_649_n 0.0394925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1175_93#_c_650_n 0.0076777f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=2.035
cc_50 VNB N_A_1175_93#_c_651_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1175_93#_c_652_n 0.0027428f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=2.405
cc_52 VNB N_A_1175_93#_c_653_n 0.00812273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1175_93#_c_654_n 0.00975764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1175_93#_c_655_n 0.00724979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1004_379#_M1007_g 0.0106845f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_56 VNB N_A_1004_379#_c_740_n 0.00699085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1004_379#_c_741_n 0.0197666f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.005
cc_58 VNB N_A_1004_379#_c_742_n 0.00621469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1004_379#_c_743_n 0.0020583f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=1.295
cc_60 VNB N_A_1004_379#_c_744_n 0.0338994f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=2.035
cc_61 VNB N_A_1004_379#_c_745_n 0.0212645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VPWR_c_814_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_432_119#_c_914_n 0.00162137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_432_119#_c_915_n 0.00633291f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_65 VNB N_A_432_119#_c_916_n 0.00252907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB Q 0.00740814f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.72
cc_67 VNB N_VGND_c_961_n 0.0109343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_962_n 0.0209936f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.005
cc_69 VNB N_VGND_c_963_n 0.00718731f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_70 VNB N_VGND_c_964_n 0.0130433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_965_n 0.0201331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_966_n 0.0126224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_967_n 0.017422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_968_n 0.0353831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_969_n 0.00372873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_970_n 0.0749189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_971_n 0.0457868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_972_n 0.0226188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_973_n 0.0172324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_974_n 0.0100021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_975_n 0.00538573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_976_n 0.459825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VPB N_CLK_M1021_g 0.0634589f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.72
cc_84 VPB CLK 0.0354669f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_85 VPB N_D_M1010_g 0.0342136f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.51
cc_86 VPB N_D_c_183_n 0.0207221f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_87 VPB N_A_240_443#_M1022_g 0.0184366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_240_443#_c_225_n 0.0146216f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_240_443#_c_235_n 0.0209062f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.005
cc_90 VPB N_A_240_443#_c_236_n 0.025234f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_91 VPB N_A_240_443#_c_227_n 0.00239476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_240_443#_c_238_n 0.00442705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_240_443#_c_239_n 0.0208439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_240_443#_c_240_n 0.00205326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_240_443#_c_241_n 0.0078704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_240_443#_c_242_n 0.0023355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_240_443#_c_228_n 0.00231488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_240_443#_c_229_n 0.0182292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_240_443#_c_245_n 0.0156045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_240_443#_c_246_n 8.42614e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_240_443#_c_231_n 0.00267824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_240_443#_c_248_n 0.00359051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_240_443#_c_249_n 9.76373e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_240_443#_c_232_n 0.0110312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_679_93#_M1005_g 0.0384892f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_106 VPB N_A_679_93#_c_386_n 0.00338499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_679_93#_c_391_n 0.00261134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_679_93#_c_392_n 0.00341104f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.005
cc_109 VPB N_A_679_93#_c_387_n 0.00483972f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.84
cc_110 VPB N_A_679_93#_c_388_n 0.0188621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_551_119#_M1011_g 0.0240555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_551_119#_c_449_n 0.0113969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_551_119#_c_452_n 0.0019585f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.005
cc_114 VPB N_A_551_119#_c_453_n 0.00870067f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.005
cc_115 VPB N_A_110_62#_M1013_g 0.0511111f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_116 VPB N_A_110_62#_c_528_n 0.125552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_110_62#_c_529_n 0.0126405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_110_62#_M1002_g 0.0434228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_110_62#_c_531_n 0.108498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_110_62#_M1014_g 0.0427155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_110_62#_c_533_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_110_62#_c_525_n 0.0272794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_110_62#_c_526_n 0.0277717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_1175_93#_c_644_n 0.00944446f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_125 VPB N_A_1175_93#_M1020_g 0.0213766f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_126 VPB N_A_1175_93#_M1008_g 0.0228149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_1175_93#_M1019_g 0.0272176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_1175_93#_c_649_n 0.0192732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_1175_93#_c_650_n 6.61225e-19 $X=-0.19 $Y=1.655 $X2=0.255
+ $Y2=2.035
cc_130 VPB N_A_1175_93#_c_652_n 0.00415381f $X=-0.19 $Y=1.655 $X2=0.255
+ $Y2=2.405
cc_131 VPB N_A_1175_93#_c_663_n 0.0193575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_1175_93#_c_664_n 0.00181377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_1175_93#_c_655_n 0.00170491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_1004_379#_M1007_g 0.0271132f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_135 VPB N_A_1004_379#_c_747_n 0.00193853f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_136 VPB N_A_1004_379#_c_748_n 0.0115258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_1004_379#_c_742_n 0.00155396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_815_n 0.0107568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_816_n 0.0206877f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.005
cc_140 VPB N_VPWR_c_817_n 0.00833896f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_141 VPB N_VPWR_c_818_n 0.00986627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_819_n 0.0384422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_820_n 0.0255792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_821_n 0.0125965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_822_n 0.00917236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_823_n 0.0560065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_824_n 0.00728331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_825_n 0.0300124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_826_n 0.0516965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_827_n 0.023482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_828_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_829_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_830_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_831_n 0.00535984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_814_n 0.110996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_432_119#_c_915_n 0.0105943f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_157 VPB Q 0.00478086f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.72
cc_158 N_CLK_c_158_n N_A_110_62#_c_515_n 0.0169316f $X=0.352 $Y=1.313 $X2=0
+ $Y2=0
cc_159 CLK N_A_110_62#_c_515_n 4.98363e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_160 CLK N_A_110_62#_c_525_n 0.129943f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_161 N_CLK_c_163_n N_A_110_62#_c_525_n 0.0331751f $X=0.352 $Y=0.84 $X2=0 $Y2=0
cc_162 N_CLK_c_160_n N_A_110_62#_c_526_n 0.0169316f $X=0.352 $Y=1.51 $X2=0 $Y2=0
cc_163 CLK N_VPWR_M1021_s 0.00269395f $X=0.155 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_164 N_CLK_M1021_g N_VPWR_c_816_n 0.0121421f $X=0.475 $Y=2.72 $X2=0 $Y2=0
cc_165 CLK N_VPWR_c_816_n 0.0238082f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_166 N_CLK_M1021_g N_VPWR_c_825_n 0.00441152f $X=0.475 $Y=2.72 $X2=0 $Y2=0
cc_167 N_CLK_M1021_g N_VPWR_c_814_n 0.00892199f $X=0.475 $Y=2.72 $X2=0 $Y2=0
cc_168 CLK N_VPWR_c_814_n 0.0015796f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_169 CLK N_VGND_c_962_n 0.0256448f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_170 N_CLK_c_162_n N_VGND_c_962_n 0.00174534f $X=0.32 $Y=1.005 $X2=0 $Y2=0
cc_171 N_CLK_c_163_n N_VGND_c_962_n 0.012443f $X=0.352 $Y=0.84 $X2=0 $Y2=0
cc_172 N_CLK_c_163_n N_VGND_c_968_n 0.00425877f $X=0.352 $Y=0.84 $X2=0 $Y2=0
cc_173 CLK N_VGND_c_976_n 0.00149307f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_174 N_CLK_c_163_n N_VGND_c_976_n 0.00861707f $X=0.352 $Y=0.84 $X2=0 $Y2=0
cc_175 N_D_c_183_n N_A_240_443#_M1004_g 0.00276112f $X=2.105 $Y=1.295 $X2=0
+ $Y2=0
cc_176 N_D_c_183_n N_A_240_443#_c_226_n 0.019256f $X=2.105 $Y=1.295 $X2=0 $Y2=0
cc_177 N_D_M1010_g N_A_240_443#_c_236_n 0.019256f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_178 N_D_M1010_g N_A_240_443#_c_227_n 6.23232e-19 $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_179 D N_A_240_443#_c_227_n 0.0261899f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_180 N_D_c_183_n N_A_240_443#_c_227_n 0.00257472f $X=2.105 $Y=1.295 $X2=0
+ $Y2=0
cc_181 N_D_c_184_n N_A_240_443#_c_227_n 6.85845e-19 $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_182 N_D_M1010_g N_A_240_443#_c_239_n 0.00544699f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_183 D N_A_240_443#_c_239_n 0.0275424f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_184 N_D_c_183_n N_A_240_443#_c_239_n 0.00846508f $X=2.105 $Y=1.295 $X2=0
+ $Y2=0
cc_185 N_D_M1010_g N_A_240_443#_c_240_n 0.0166295f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_186 N_D_M1010_g N_A_240_443#_c_241_n 0.00664286f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_187 N_D_M1010_g N_A_240_443#_c_242_n 2.84307e-19 $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_188 N_D_M1010_g N_A_240_443#_c_228_n 7.82885e-19 $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_189 N_D_M1010_g N_A_110_62#_M1013_g 0.00944498f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_190 D N_A_110_62#_M1013_g 0.00136203f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_191 N_D_c_183_n N_A_110_62#_M1013_g 0.0148551f $X=2.105 $Y=1.295 $X2=0 $Y2=0
cc_192 D N_A_110_62#_M1009_g 9.65644e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_193 N_D_c_183_n N_A_110_62#_M1009_g 0.01631f $X=2.105 $Y=1.295 $X2=0 $Y2=0
cc_194 N_D_c_184_n N_A_110_62#_M1009_g 0.0117234f $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_195 N_D_M1010_g N_A_110_62#_c_528_n 0.00532498f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_196 N_D_c_184_n N_A_110_62#_c_518_n 0.0103107f $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_197 N_D_c_183_n N_A_110_62#_M1015_g 9.4343e-19 $X=2.105 $Y=1.295 $X2=0 $Y2=0
cc_198 N_D_c_184_n N_A_110_62#_M1015_g 0.0151193f $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_199 N_D_M1010_g N_VPWR_c_817_n 0.00146359f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_200 N_D_M1010_g N_A_432_119#_c_914_n 0.00655307f $X=2.32 $Y=2.425 $X2=0 $Y2=0
cc_201 D N_A_432_119#_c_919_n 0.00360215f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_202 N_D_c_183_n N_A_432_119#_c_919_n 0.00683183f $X=2.105 $Y=1.295 $X2=0
+ $Y2=0
cc_203 N_D_c_184_n N_A_432_119#_c_919_n 0.00320787f $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_204 D N_A_432_119#_c_916_n 0.047266f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_205 N_D_c_183_n N_A_432_119#_c_916_n 0.00655307f $X=2.105 $Y=1.295 $X2=0
+ $Y2=0
cc_206 N_D_c_184_n N_A_432_119#_c_916_n 0.00314603f $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_207 D N_VGND_c_963_n 0.0054005f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_208 N_D_c_183_n N_VGND_c_963_n 0.00174559f $X=2.105 $Y=1.295 $X2=0 $Y2=0
cc_209 N_D_c_184_n N_VGND_c_963_n 0.00909379f $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_210 N_D_c_184_n N_VGND_c_976_n 7.88961e-19 $X=2.167 $Y=1.13 $X2=0 $Y2=0
cc_211 N_A_240_443#_c_265_p N_A_679_93#_M1011_d 0.00746136f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_212 N_A_240_443#_M1004_g N_A_679_93#_M1024_g 0.0321048f $X=3.11 $Y=0.805
+ $X2=0 $Y2=0
cc_213 N_A_240_443#_c_229_n N_A_679_93#_M1005_g 0.00317137f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_214 N_A_240_443#_c_246_n N_A_679_93#_M1005_g 0.00156732f $X=3.605 $Y=2.76
+ $X2=0 $Y2=0
cc_215 N_A_240_443#_c_265_p N_A_679_93#_M1005_g 0.0116167f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_216 N_A_240_443#_c_265_p N_A_679_93#_c_391_n 0.0391313f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_217 N_A_240_443#_c_265_p N_A_679_93#_c_392_n 0.0159285f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_218 N_A_240_443#_c_272_p N_A_679_93#_c_392_n 0.00728045f $X=3.69 $Y=2.37
+ $X2=0 $Y2=0
cc_219 N_A_240_443#_c_265_p N_A_679_93#_c_403_n 0.0176317f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_220 N_A_240_443#_M1018_g N_A_679_93#_c_387_n 0.0119637f $X=5.02 $Y=0.805
+ $X2=0 $Y2=0
cc_221 N_A_240_443#_c_230_n N_A_679_93#_c_387_n 0.0196832f $X=5.075 $Y=1.555
+ $X2=0 $Y2=0
cc_222 N_A_240_443#_c_231_n N_A_679_93#_c_387_n 0.0258981f $X=5.075 $Y=2.285
+ $X2=0 $Y2=0
cc_223 N_A_240_443#_c_226_n N_A_679_93#_c_388_n 0.0321048f $X=2.93 $Y=1.535
+ $X2=0 $Y2=0
cc_224 N_A_240_443#_c_229_n N_A_679_93#_c_388_n 0.0060803f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_225 N_A_240_443#_c_272_p N_A_679_93#_c_388_n 0.00183179f $X=3.69 $Y=2.37
+ $X2=0 $Y2=0
cc_226 N_A_240_443#_c_228_n N_A_551_119#_M1022_d 0.00407654f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_227 N_A_240_443#_c_265_p N_A_551_119#_M1011_g 0.0125701f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_228 N_A_240_443#_c_231_n N_A_551_119#_M1011_g 5.77305e-19 $X=5.075 $Y=2.285
+ $X2=0 $Y2=0
cc_229 N_A_240_443#_M1022_g N_A_551_119#_c_449_n 0.00156175f $X=2.75 $Y=2.425
+ $X2=0 $Y2=0
cc_230 N_A_240_443#_M1004_g N_A_551_119#_c_449_n 0.00418913f $X=3.11 $Y=0.805
+ $X2=0 $Y2=0
cc_231 N_A_240_443#_c_226_n N_A_551_119#_c_449_n 0.00469832f $X=2.93 $Y=1.535
+ $X2=0 $Y2=0
cc_232 N_A_240_443#_c_228_n N_A_551_119#_c_449_n 0.0880137f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_233 N_A_240_443#_c_229_n N_A_551_119#_c_449_n 0.00576972f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_234 N_A_240_443#_c_245_n N_A_551_119#_c_449_n 0.0153109f $X=3.52 $Y=2.85
+ $X2=0 $Y2=0
cc_235 N_A_240_443#_M1004_g N_A_551_119#_c_451_n 0.0189802f $X=3.11 $Y=0.805
+ $X2=0 $Y2=0
cc_236 N_A_240_443#_c_226_n N_A_551_119#_c_451_n 0.00397144f $X=2.93 $Y=1.535
+ $X2=0 $Y2=0
cc_237 N_A_240_443#_c_228_n N_A_551_119#_c_451_n 0.00834417f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_238 N_A_240_443#_c_232_n N_A_551_119#_c_453_n 0.0111415f $X=5.14 $Y=1.39
+ $X2=0 $Y2=0
cc_239 N_A_240_443#_M1018_g N_A_551_119#_c_454_n 0.0100286f $X=5.02 $Y=0.805
+ $X2=0 $Y2=0
cc_240 N_A_240_443#_c_227_n N_A_110_62#_c_514_n 0.0154655f $X=1.42 $Y=0.805
+ $X2=0 $Y2=0
cc_241 N_A_240_443#_c_227_n N_A_110_62#_M1013_g 0.0193828f $X=1.42 $Y=0.805
+ $X2=0 $Y2=0
cc_242 N_A_240_443#_c_238_n N_A_110_62#_M1013_g 0.00337022f $X=1.325 $Y=2.36
+ $X2=0 $Y2=0
cc_243 N_A_240_443#_c_239_n N_A_110_62#_M1013_g 0.00561898f $X=2.09 $Y=2.02
+ $X2=0 $Y2=0
cc_244 N_A_240_443#_c_240_n N_A_110_62#_M1013_g 0.00119138f $X=2.18 $Y=2.76
+ $X2=0 $Y2=0
cc_245 N_A_240_443#_c_242_n N_A_110_62#_M1013_g 5.18129e-19 $X=2.27 $Y=2.85
+ $X2=0 $Y2=0
cc_246 N_A_240_443#_c_248_n N_A_110_62#_M1013_g 0.0113953f $X=1.397 $Y=2.02
+ $X2=0 $Y2=0
cc_247 N_A_240_443#_c_227_n N_A_110_62#_M1009_g 0.0117219f $X=1.42 $Y=0.805
+ $X2=0 $Y2=0
cc_248 N_A_240_443#_M1022_g N_A_110_62#_c_528_n 0.00532498f $X=2.75 $Y=2.425
+ $X2=0 $Y2=0
cc_249 N_A_240_443#_c_241_n N_A_110_62#_c_528_n 0.00802429f $X=2.8 $Y=2.85 $X2=0
+ $Y2=0
cc_250 N_A_240_443#_c_242_n N_A_110_62#_c_528_n 0.00381984f $X=2.27 $Y=2.85
+ $X2=0 $Y2=0
cc_251 N_A_240_443#_c_245_n N_A_110_62#_c_528_n 0.00679584f $X=3.52 $Y=2.85
+ $X2=0 $Y2=0
cc_252 N_A_240_443#_c_249_n N_A_110_62#_c_528_n 0.00358867f $X=2.885 $Y=2.85
+ $X2=0 $Y2=0
cc_253 N_A_240_443#_M1004_g N_A_110_62#_M1015_g 0.0131996f $X=3.11 $Y=0.805
+ $X2=0 $Y2=0
cc_254 N_A_240_443#_c_226_n N_A_110_62#_M1015_g 0.00592368f $X=2.93 $Y=1.535
+ $X2=0 $Y2=0
cc_255 N_A_240_443#_M1004_g N_A_110_62#_c_521_n 0.0100275f $X=3.11 $Y=0.805
+ $X2=0 $Y2=0
cc_256 N_A_240_443#_M1018_g N_A_110_62#_c_521_n 0.0104164f $X=5.02 $Y=0.805
+ $X2=0 $Y2=0
cc_257 N_A_240_443#_M1022_g N_A_110_62#_M1002_g 0.00747449f $X=2.75 $Y=2.425
+ $X2=0 $Y2=0
cc_258 N_A_240_443#_c_228_n N_A_110_62#_M1002_g 0.00193823f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_259 N_A_240_443#_c_245_n N_A_110_62#_M1002_g 0.0181028f $X=3.52 $Y=2.85 $X2=0
+ $Y2=0
cc_260 N_A_240_443#_c_246_n N_A_110_62#_M1002_g 0.00601997f $X=3.605 $Y=2.76
+ $X2=0 $Y2=0
cc_261 N_A_240_443#_c_272_p N_A_110_62#_M1002_g 0.00318855f $X=3.69 $Y=2.37
+ $X2=0 $Y2=0
cc_262 N_A_240_443#_c_245_n N_A_110_62#_c_531_n 0.00172486f $X=3.52 $Y=2.85
+ $X2=0 $Y2=0
cc_263 N_A_240_443#_c_265_p N_A_110_62#_c_531_n 0.00844611f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_264 N_A_240_443#_c_235_n N_A_110_62#_M1014_g 0.00688796f $X=5.74 $Y=1.785
+ $X2=0 $Y2=0
cc_265 N_A_240_443#_c_265_p N_A_110_62#_M1014_g 0.018642f $X=4.985 $Y=2.37 $X2=0
+ $Y2=0
cc_266 N_A_240_443#_c_231_n N_A_110_62#_M1014_g 0.0141726f $X=5.075 $Y=2.285
+ $X2=0 $Y2=0
cc_267 N_A_240_443#_c_232_n N_A_110_62#_M1014_g 0.0066561f $X=5.14 $Y=1.39 $X2=0
+ $Y2=0
cc_268 N_A_240_443#_M1018_g N_A_110_62#_M1006_g 0.0175305f $X=5.02 $Y=0.805
+ $X2=0 $Y2=0
cc_269 N_A_240_443#_c_225_n N_A_110_62#_M1006_g 0.00300439f $X=5.665 $Y=1.71
+ $X2=0 $Y2=0
cc_270 N_A_240_443#_c_227_n N_A_110_62#_c_523_n 0.00619557f $X=1.42 $Y=0.805
+ $X2=0 $Y2=0
cc_271 N_A_240_443#_c_239_n N_A_110_62#_c_523_n 0.00319484f $X=2.09 $Y=2.02
+ $X2=0 $Y2=0
cc_272 N_A_240_443#_c_227_n N_A_110_62#_c_525_n 0.107787f $X=1.42 $Y=0.805 $X2=0
+ $Y2=0
cc_273 N_A_240_443#_c_238_n N_A_110_62#_c_525_n 0.0617213f $X=1.325 $Y=2.36
+ $X2=0 $Y2=0
cc_274 N_A_240_443#_c_248_n N_A_110_62#_c_525_n 0.0153667f $X=1.397 $Y=2.02
+ $X2=0 $Y2=0
cc_275 N_A_240_443#_c_227_n N_A_110_62#_c_526_n 0.00453047f $X=1.42 $Y=0.805
+ $X2=0 $Y2=0
cc_276 N_A_240_443#_c_232_n N_A_1175_93#_M1001_g 0.00252037f $X=5.14 $Y=1.39
+ $X2=0 $Y2=0
cc_277 N_A_240_443#_c_225_n N_A_1175_93#_c_644_n 0.0239425f $X=5.665 $Y=1.71
+ $X2=0 $Y2=0
cc_278 N_A_240_443#_c_232_n N_A_1175_93#_c_644_n 0.00300984f $X=5.14 $Y=1.39
+ $X2=0 $Y2=0
cc_279 N_A_240_443#_c_235_n N_A_1175_93#_M1020_g 0.0239425f $X=5.74 $Y=1.785
+ $X2=0 $Y2=0
cc_280 N_A_240_443#_c_225_n N_A_1175_93#_c_664_n 7.03886e-19 $X=5.665 $Y=1.71
+ $X2=0 $Y2=0
cc_281 N_A_240_443#_c_265_p N_A_1004_379#_M1014_d 0.00561276f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_282 N_A_240_443#_c_231_n N_A_1004_379#_M1014_d 0.00369051f $X=5.075 $Y=2.285
+ $X2=0 $Y2=0
cc_283 N_A_240_443#_c_231_n N_A_1004_379#_c_747_n 0.0313664f $X=5.075 $Y=2.285
+ $X2=0 $Y2=0
cc_284 N_A_240_443#_c_232_n N_A_1004_379#_c_747_n 0.00698611f $X=5.14 $Y=1.39
+ $X2=0 $Y2=0
cc_285 N_A_240_443#_c_265_p N_A_1004_379#_c_748_n 0.0144464f $X=4.985 $Y=2.37
+ $X2=0 $Y2=0
cc_286 N_A_240_443#_M1018_g N_A_1004_379#_c_740_n 0.00665882f $X=5.02 $Y=0.805
+ $X2=0 $Y2=0
cc_287 N_A_240_443#_c_225_n N_A_1004_379#_c_740_n 0.00203504f $X=5.665 $Y=1.71
+ $X2=0 $Y2=0
cc_288 N_A_240_443#_c_230_n N_A_1004_379#_c_740_n 0.0130747f $X=5.075 $Y=1.555
+ $X2=0 $Y2=0
cc_289 N_A_240_443#_c_232_n N_A_1004_379#_c_740_n 0.0103303f $X=5.14 $Y=1.39
+ $X2=0 $Y2=0
cc_290 N_A_240_443#_c_225_n N_A_1004_379#_c_741_n 0.00536119f $X=5.665 $Y=1.71
+ $X2=0 $Y2=0
cc_291 N_A_240_443#_c_225_n N_A_1004_379#_c_742_n 0.0136512f $X=5.665 $Y=1.71
+ $X2=0 $Y2=0
cc_292 N_A_240_443#_c_235_n N_A_1004_379#_c_742_n 0.00913853f $X=5.74 $Y=1.785
+ $X2=0 $Y2=0
cc_293 N_A_240_443#_c_230_n N_A_1004_379#_c_742_n 0.018753f $X=5.075 $Y=1.555
+ $X2=0 $Y2=0
cc_294 N_A_240_443#_c_231_n N_A_1004_379#_c_742_n 0.0149652f $X=5.075 $Y=2.285
+ $X2=0 $Y2=0
cc_295 N_A_240_443#_c_232_n N_A_1004_379#_c_742_n 0.00335117f $X=5.14 $Y=1.39
+ $X2=0 $Y2=0
cc_296 N_A_240_443#_c_240_n N_VPWR_M1013_d 0.00443199f $X=2.18 $Y=2.76 $X2=0
+ $Y2=0
cc_297 N_A_240_443#_c_265_p N_VPWR_M1005_d 0.00857734f $X=4.985 $Y=2.37 $X2=0
+ $Y2=0
cc_298 N_A_240_443#_c_238_n N_VPWR_c_817_n 0.0221126f $X=1.325 $Y=2.36 $X2=0
+ $Y2=0
cc_299 N_A_240_443#_c_239_n N_VPWR_c_817_n 0.0233644f $X=2.09 $Y=2.02 $X2=0
+ $Y2=0
cc_300 N_A_240_443#_c_240_n N_VPWR_c_817_n 0.0367701f $X=2.18 $Y=2.76 $X2=0
+ $Y2=0
cc_301 N_A_240_443#_c_242_n N_VPWR_c_817_n 0.0159229f $X=2.27 $Y=2.85 $X2=0
+ $Y2=0
cc_302 N_A_240_443#_c_245_n N_VPWR_c_818_n 0.0111029f $X=3.52 $Y=2.85 $X2=0
+ $Y2=0
cc_303 N_A_240_443#_c_246_n N_VPWR_c_818_n 0.00712924f $X=3.605 $Y=2.76 $X2=0
+ $Y2=0
cc_304 N_A_240_443#_c_265_p N_VPWR_c_818_n 0.0266042f $X=4.985 $Y=2.37 $X2=0
+ $Y2=0
cc_305 N_A_240_443#_c_235_n N_VPWR_c_819_n 0.00130302f $X=5.74 $Y=1.785 $X2=0
+ $Y2=0
cc_306 N_A_240_443#_c_238_n N_VPWR_c_825_n 0.00632433f $X=1.325 $Y=2.36 $X2=0
+ $Y2=0
cc_307 N_A_240_443#_c_241_n N_VPWR_c_826_n 0.0184625f $X=2.8 $Y=2.85 $X2=0 $Y2=0
cc_308 N_A_240_443#_c_242_n N_VPWR_c_826_n 0.00690996f $X=2.27 $Y=2.85 $X2=0
+ $Y2=0
cc_309 N_A_240_443#_c_245_n N_VPWR_c_826_n 0.0253157f $X=3.52 $Y=2.85 $X2=0
+ $Y2=0
cc_310 N_A_240_443#_c_249_n N_VPWR_c_826_n 0.00652607f $X=2.885 $Y=2.85 $X2=0
+ $Y2=0
cc_311 N_A_240_443#_c_235_n N_VPWR_c_814_n 0.00373935f $X=5.74 $Y=1.785 $X2=0
+ $Y2=0
cc_312 N_A_240_443#_c_238_n N_VPWR_c_814_n 0.00713006f $X=1.325 $Y=2.36 $X2=0
+ $Y2=0
cc_313 N_A_240_443#_c_241_n N_VPWR_c_814_n 0.0161173f $X=2.8 $Y=2.85 $X2=0 $Y2=0
cc_314 N_A_240_443#_c_242_n N_VPWR_c_814_n 0.00576321f $X=2.27 $Y=2.85 $X2=0
+ $Y2=0
cc_315 N_A_240_443#_c_245_n N_VPWR_c_814_n 0.0219808f $X=3.52 $Y=2.85 $X2=0
+ $Y2=0
cc_316 N_A_240_443#_c_249_n N_VPWR_c_814_n 0.00544303f $X=2.885 $Y=2.85 $X2=0
+ $Y2=0
cc_317 N_A_240_443#_M1004_g N_A_432_119#_c_914_n 0.00136126f $X=3.11 $Y=0.805
+ $X2=0 $Y2=0
cc_318 N_A_240_443#_c_226_n N_A_432_119#_c_915_n 0.00675711f $X=2.93 $Y=1.535
+ $X2=0 $Y2=0
cc_319 N_A_240_443#_c_239_n N_A_432_119#_c_915_n 0.0136934f $X=2.09 $Y=2.02
+ $X2=0 $Y2=0
cc_320 N_A_240_443#_c_240_n N_A_432_119#_c_915_n 0.0207187f $X=2.18 $Y=2.76
+ $X2=0 $Y2=0
cc_321 N_A_240_443#_c_241_n N_A_432_119#_c_915_n 0.0140896f $X=2.8 $Y=2.85 $X2=0
+ $Y2=0
cc_322 N_A_240_443#_c_228_n N_A_432_119#_c_915_n 0.0724579f $X=2.885 $Y=1.55
+ $X2=0 $Y2=0
cc_323 N_A_240_443#_M1004_g N_A_432_119#_c_916_n 9.59776e-19 $X=3.11 $Y=0.805
+ $X2=0 $Y2=0
cc_324 N_A_240_443#_c_272_p A_705_443# 0.00115303f $X=3.69 $Y=2.37 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A_240_443#_c_227_n N_VGND_c_968_n 0.0066463f $X=1.42 $Y=0.805 $X2=0
+ $Y2=0
cc_326 N_A_240_443#_M1004_g N_VGND_c_970_n 0.00149099f $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_327 N_A_240_443#_M1018_g N_VGND_c_970_n 5.98494e-19 $X=5.02 $Y=0.805 $X2=0
+ $Y2=0
cc_328 N_A_240_443#_M1004_g N_VGND_c_976_n 9.39239e-19 $X=3.11 $Y=0.805 $X2=0
+ $Y2=0
cc_329 N_A_240_443#_M1018_g N_VGND_c_976_n 9.39239e-19 $X=5.02 $Y=0.805 $X2=0
+ $Y2=0
cc_330 N_A_240_443#_c_227_n N_VGND_c_976_n 0.0112435f $X=1.42 $Y=0.805 $X2=0
+ $Y2=0
cc_331 N_A_679_93#_M1005_g N_A_551_119#_M1011_g 0.0235527f $X=3.81 $Y=2.425
+ $X2=0 $Y2=0
cc_332 N_A_679_93#_c_386_n N_A_551_119#_M1011_g 0.00177413f $X=3.77 $Y=1.57
+ $X2=0 $Y2=0
cc_333 N_A_679_93#_c_391_n N_A_551_119#_M1011_g 0.0130978f $X=4.595 $Y=2.015
+ $X2=0 $Y2=0
cc_334 N_A_679_93#_c_387_n N_A_551_119#_M1011_g 0.00435735f $X=4.71 $Y=0.75
+ $X2=0 $Y2=0
cc_335 N_A_679_93#_c_388_n N_A_551_119#_M1011_g 0.00162817f $X=3.81 $Y=1.57
+ $X2=0 $Y2=0
cc_336 N_A_679_93#_M1024_g N_A_551_119#_c_449_n 0.00770366f $X=3.47 $Y=0.805
+ $X2=0 $Y2=0
cc_337 N_A_679_93#_M1005_g N_A_551_119#_c_449_n 0.00121054f $X=3.81 $Y=2.425
+ $X2=0 $Y2=0
cc_338 N_A_679_93#_c_386_n N_A_551_119#_c_449_n 0.0295082f $X=3.77 $Y=1.57 $X2=0
+ $Y2=0
cc_339 N_A_679_93#_c_392_n N_A_551_119#_c_449_n 0.0128999f $X=3.935 $Y=2.015
+ $X2=0 $Y2=0
cc_340 N_A_679_93#_M1024_g N_A_551_119#_c_450_n 0.0198717f $X=3.47 $Y=0.805
+ $X2=0 $Y2=0
cc_341 N_A_679_93#_c_386_n N_A_551_119#_c_450_n 0.0251839f $X=3.77 $Y=1.57 $X2=0
+ $Y2=0
cc_342 N_A_679_93#_c_388_n N_A_551_119#_c_450_n 0.00453691f $X=3.81 $Y=1.57
+ $X2=0 $Y2=0
cc_343 N_A_679_93#_M1024_g N_A_551_119#_c_451_n 0.00213312f $X=3.47 $Y=0.805
+ $X2=0 $Y2=0
cc_344 N_A_679_93#_M1024_g N_A_551_119#_c_452_n 0.00295111f $X=3.47 $Y=0.805
+ $X2=0 $Y2=0
cc_345 N_A_679_93#_c_386_n N_A_551_119#_c_452_n 0.0150617f $X=3.77 $Y=1.57 $X2=0
+ $Y2=0
cc_346 N_A_679_93#_c_391_n N_A_551_119#_c_452_n 0.0131786f $X=4.595 $Y=2.015
+ $X2=0 $Y2=0
cc_347 N_A_679_93#_c_387_n N_A_551_119#_c_452_n 0.0331652f $X=4.71 $Y=0.75 $X2=0
+ $Y2=0
cc_348 N_A_679_93#_c_388_n N_A_551_119#_c_452_n 0.00109276f $X=3.81 $Y=1.57
+ $X2=0 $Y2=0
cc_349 N_A_679_93#_M1024_g N_A_551_119#_c_453_n 0.00125981f $X=3.47 $Y=0.805
+ $X2=0 $Y2=0
cc_350 N_A_679_93#_c_386_n N_A_551_119#_c_453_n 0.00102834f $X=3.77 $Y=1.57
+ $X2=0 $Y2=0
cc_351 N_A_679_93#_c_391_n N_A_551_119#_c_453_n 0.00246492f $X=4.595 $Y=2.015
+ $X2=0 $Y2=0
cc_352 N_A_679_93#_c_388_n N_A_551_119#_c_453_n 0.0147099f $X=3.81 $Y=1.57 $X2=0
+ $Y2=0
cc_353 N_A_679_93#_c_387_n N_A_551_119#_c_454_n 0.00497528f $X=4.71 $Y=0.75
+ $X2=0 $Y2=0
cc_354 N_A_679_93#_M1024_g N_A_110_62#_c_521_n 0.0103107f $X=3.47 $Y=0.805 $X2=0
+ $Y2=0
cc_355 N_A_679_93#_c_387_n N_A_110_62#_c_521_n 0.00419295f $X=4.71 $Y=0.75 $X2=0
+ $Y2=0
cc_356 N_A_679_93#_M1005_g N_A_110_62#_M1002_g 0.0412126f $X=3.81 $Y=2.425 $X2=0
+ $Y2=0
cc_357 N_A_679_93#_c_392_n N_A_110_62#_M1002_g 2.51516e-19 $X=3.935 $Y=2.015
+ $X2=0 $Y2=0
cc_358 N_A_679_93#_c_388_n N_A_110_62#_M1002_g 0.00681352f $X=3.81 $Y=1.57 $X2=0
+ $Y2=0
cc_359 N_A_679_93#_M1005_g N_A_110_62#_c_531_n 0.00640451f $X=3.81 $Y=2.425
+ $X2=0 $Y2=0
cc_360 N_A_679_93#_c_387_n N_A_110_62#_M1014_g 0.00121736f $X=4.71 $Y=0.75 $X2=0
+ $Y2=0
cc_361 N_A_679_93#_c_387_n N_A_1004_379#_c_740_n 0.0138223f $X=4.71 $Y=0.75
+ $X2=0 $Y2=0
cc_362 N_A_679_93#_c_391_n N_VPWR_M1005_d 0.0128577f $X=4.595 $Y=2.015 $X2=0
+ $Y2=0
cc_363 N_A_679_93#_M1005_g N_VPWR_c_818_n 0.00152978f $X=3.81 $Y=2.425 $X2=0
+ $Y2=0
cc_364 N_A_679_93#_M1005_g N_VPWR_c_814_n 9.66522e-19 $X=3.81 $Y=2.425 $X2=0
+ $Y2=0
cc_365 N_A_679_93#_M1024_g N_VGND_c_970_n 0.0107156f $X=3.47 $Y=0.805 $X2=0
+ $Y2=0
cc_366 N_A_679_93#_c_387_n N_VGND_c_970_n 0.0129272f $X=4.71 $Y=0.75 $X2=0 $Y2=0
cc_367 N_A_679_93#_c_387_n N_VGND_c_971_n 0.00468217f $X=4.71 $Y=0.75 $X2=0
+ $Y2=0
cc_368 N_A_679_93#_M1024_g N_VGND_c_976_n 7.88961e-19 $X=3.47 $Y=0.805 $X2=0
+ $Y2=0
cc_369 N_A_679_93#_c_387_n N_VGND_c_976_n 0.00572408f $X=4.71 $Y=0.75 $X2=0
+ $Y2=0
cc_370 N_A_551_119#_c_451_n N_A_110_62#_M1015_g 5.60804e-19 $X=3.35 $Y=1.14
+ $X2=0 $Y2=0
cc_371 N_A_551_119#_c_451_n N_A_110_62#_c_521_n 0.00681752f $X=3.35 $Y=1.14
+ $X2=0 $Y2=0
cc_372 N_A_551_119#_c_454_n N_A_110_62#_c_521_n 0.0104018f $X=4.372 $Y=1.345
+ $X2=0 $Y2=0
cc_373 N_A_551_119#_c_449_n N_A_110_62#_M1002_g 0.00338226f $X=3.235 $Y=2.425
+ $X2=0 $Y2=0
cc_374 N_A_551_119#_M1011_g N_A_110_62#_c_531_n 0.0100858f $X=4.435 $Y=2.315
+ $X2=0 $Y2=0
cc_375 N_A_551_119#_M1011_g N_A_110_62#_M1014_g 0.0312813f $X=4.435 $Y=2.315
+ $X2=0 $Y2=0
cc_376 N_A_551_119#_M1011_g N_VPWR_c_818_n 0.00579056f $X=4.435 $Y=2.315 $X2=0
+ $Y2=0
cc_377 N_A_551_119#_M1011_g N_VPWR_c_814_n 9.39239e-19 $X=4.435 $Y=2.315 $X2=0
+ $Y2=0
cc_378 N_A_551_119#_c_449_n N_A_432_119#_c_914_n 0.00509621f $X=3.235 $Y=2.425
+ $X2=0 $Y2=0
cc_379 N_A_551_119#_c_451_n N_A_432_119#_c_916_n 0.00895227f $X=3.35 $Y=1.14
+ $X2=0 $Y2=0
cc_380 N_A_551_119#_c_450_n N_VGND_M1024_d 0.00459726f $X=4.175 $Y=1.14 $X2=0
+ $Y2=0
cc_381 N_A_551_119#_c_450_n N_VGND_c_970_n 0.0683622f $X=4.175 $Y=1.14 $X2=0
+ $Y2=0
cc_382 N_A_551_119#_c_451_n N_VGND_c_970_n 0.0121023f $X=3.35 $Y=1.14 $X2=0
+ $Y2=0
cc_383 N_A_551_119#_c_453_n N_VGND_c_970_n 9.25537e-19 $X=4.34 $Y=1.51 $X2=0
+ $Y2=0
cc_384 N_A_551_119#_c_454_n N_VGND_c_970_n 0.00815768f $X=4.372 $Y=1.345 $X2=0
+ $Y2=0
cc_385 N_A_551_119#_c_451_n N_VGND_c_976_n 0.0157494f $X=3.35 $Y=1.14 $X2=0
+ $Y2=0
cc_386 N_A_551_119#_c_454_n N_VGND_c_976_n 9.14192e-19 $X=4.372 $Y=1.345 $X2=0
+ $Y2=0
cc_387 N_A_551_119#_c_451_n A_637_119# 0.00103048f $X=3.35 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A_110_62#_M1006_g N_A_1175_93#_M1001_g 0.0397709f $X=5.59 $Y=0.805
+ $X2=0 $Y2=0
cc_389 N_A_110_62#_M1014_g N_A_1004_379#_c_747_n 0.0018309f $X=4.945 $Y=2.315
+ $X2=0 $Y2=0
cc_390 N_A_110_62#_M1014_g N_A_1004_379#_c_748_n 0.009497f $X=4.945 $Y=2.315
+ $X2=0 $Y2=0
cc_391 N_A_110_62#_c_521_n N_A_1004_379#_c_740_n 0.00520438f $X=5.515 $Y=0.18
+ $X2=0 $Y2=0
cc_392 N_A_110_62#_M1006_g N_A_1004_379#_c_740_n 0.0242914f $X=5.59 $Y=0.805
+ $X2=0 $Y2=0
cc_393 N_A_110_62#_M1006_g N_A_1004_379#_c_741_n 6.70695e-19 $X=5.59 $Y=0.805
+ $X2=0 $Y2=0
cc_394 N_A_110_62#_M1014_g N_A_1004_379#_c_742_n 2.89935e-19 $X=4.945 $Y=2.315
+ $X2=0 $Y2=0
cc_395 N_A_110_62#_c_525_n N_VPWR_c_816_n 0.0150255f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_396 N_A_110_62#_M1013_g N_VPWR_c_817_n 0.0156675f $X=1.54 $Y=2.535 $X2=0
+ $Y2=0
cc_397 N_A_110_62#_c_528_n N_VPWR_c_817_n 0.0187754f $X=3.375 $Y=3.15 $X2=0
+ $Y2=0
cc_398 N_A_110_62#_c_529_n N_VPWR_c_817_n 0.00388727f $X=1.615 $Y=3.15 $X2=0
+ $Y2=0
cc_399 N_A_110_62#_c_525_n N_VPWR_c_817_n 0.00620939f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_400 N_A_110_62#_M1002_g N_VPWR_c_818_n 0.00463142f $X=3.45 $Y=2.425 $X2=0
+ $Y2=0
cc_401 N_A_110_62#_c_531_n N_VPWR_c_818_n 0.0254884f $X=4.87 $Y=3.15 $X2=0 $Y2=0
cc_402 N_A_110_62#_M1014_g N_VPWR_c_818_n 0.00564751f $X=4.945 $Y=2.315 $X2=0
+ $Y2=0
cc_403 N_A_110_62#_c_531_n N_VPWR_c_823_n 0.026094f $X=4.87 $Y=3.15 $X2=0 $Y2=0
cc_404 N_A_110_62#_c_529_n N_VPWR_c_825_n 0.00486043f $X=1.615 $Y=3.15 $X2=0
+ $Y2=0
cc_405 N_A_110_62#_c_525_n N_VPWR_c_825_n 0.0274154f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_406 N_A_110_62#_c_528_n N_VPWR_c_826_n 0.0522558f $X=3.375 $Y=3.15 $X2=0
+ $Y2=0
cc_407 N_A_110_62#_c_528_n N_VPWR_c_814_n 0.0398638f $X=3.375 $Y=3.15 $X2=0
+ $Y2=0
cc_408 N_A_110_62#_c_529_n N_VPWR_c_814_n 0.00983503f $X=1.615 $Y=3.15 $X2=0
+ $Y2=0
cc_409 N_A_110_62#_c_531_n N_VPWR_c_814_n 0.0556786f $X=4.87 $Y=3.15 $X2=0 $Y2=0
cc_410 N_A_110_62#_c_533_n N_VPWR_c_814_n 0.00381437f $X=3.45 $Y=3.15 $X2=0
+ $Y2=0
cc_411 N_A_110_62#_c_525_n N_VPWR_c_814_n 0.0170136f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_412 N_A_110_62#_M1015_g N_A_432_119#_c_914_n 4.82938e-19 $X=2.68 $Y=0.805
+ $X2=0 $Y2=0
cc_413 N_A_110_62#_c_518_n N_A_432_119#_c_919_n 0.00531785f $X=2.605 $Y=0.18
+ $X2=0 $Y2=0
cc_414 N_A_110_62#_M1015_g N_A_432_119#_c_919_n 0.00837958f $X=2.68 $Y=0.805
+ $X2=0 $Y2=0
cc_415 N_A_110_62#_M1015_g N_A_432_119#_c_916_n 0.00470141f $X=2.68 $Y=0.805
+ $X2=0 $Y2=0
cc_416 N_A_110_62#_M1009_g N_VGND_c_963_n 0.0125142f $X=1.655 $Y=0.805 $X2=0
+ $Y2=0
cc_417 N_A_110_62#_c_518_n N_VGND_c_963_n 0.0207766f $X=2.605 $Y=0.18 $X2=0
+ $Y2=0
cc_418 N_A_110_62#_M1015_g N_VGND_c_963_n 0.00603465f $X=2.68 $Y=0.805 $X2=0
+ $Y2=0
cc_419 N_A_110_62#_c_521_n N_VGND_c_964_n 0.0106506f $X=5.515 $Y=0.18 $X2=0
+ $Y2=0
cc_420 N_A_110_62#_M1006_g N_VGND_c_964_n 0.00165446f $X=5.59 $Y=0.805 $X2=0
+ $Y2=0
cc_421 N_A_110_62#_c_519_n N_VGND_c_968_n 0.00674787f $X=1.73 $Y=0.18 $X2=0
+ $Y2=0
cc_422 N_A_110_62#_c_525_n N_VGND_c_968_n 0.0209697f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_423 N_A_110_62#_c_518_n N_VGND_c_970_n 0.046512f $X=2.605 $Y=0.18 $X2=0 $Y2=0
cc_424 N_A_110_62#_c_521_n N_VGND_c_970_n 0.0576204f $X=5.515 $Y=0.18 $X2=0
+ $Y2=0
cc_425 N_A_110_62#_c_521_n N_VGND_c_971_n 0.0369091f $X=5.515 $Y=0.18 $X2=0
+ $Y2=0
cc_426 N_A_110_62#_c_518_n N_VGND_c_976_n 0.0191747f $X=2.605 $Y=0.18 $X2=0
+ $Y2=0
cc_427 N_A_110_62#_c_519_n N_VGND_c_976_n 0.0112172f $X=1.73 $Y=0.18 $X2=0 $Y2=0
cc_428 N_A_110_62#_c_521_n N_VGND_c_976_n 0.0683789f $X=5.515 $Y=0.18 $X2=0
+ $Y2=0
cc_429 N_A_110_62#_c_524_n N_VGND_c_976_n 0.00877294f $X=2.68 $Y=0.18 $X2=0
+ $Y2=0
cc_430 N_A_110_62#_c_525_n N_VGND_c_976_n 0.0165556f $X=0.69 $Y=0.495 $X2=0
+ $Y2=0
cc_431 N_A_1175_93#_M1020_g N_A_1004_379#_M1007_g 0.0135165f $X=6.1 $Y=2.105
+ $X2=0 $Y2=0
cc_432 N_A_1175_93#_c_649_n N_A_1004_379#_M1007_g 0.00590454f $X=7.63 $Y=1.51
+ $X2=0 $Y2=0
cc_433 N_A_1175_93#_c_652_n N_A_1004_379#_M1007_g 0.0162042f $X=6.75 $Y=1.72
+ $X2=0 $Y2=0
cc_434 N_A_1175_93#_c_663_n N_A_1004_379#_M1007_g 0.00754364f $X=6.855 $Y=2.04
+ $X2=0 $Y2=0
cc_435 N_A_1175_93#_c_664_n N_A_1004_379#_M1007_g 8.38198e-19 $X=6.19 $Y=1.56
+ $X2=0 $Y2=0
cc_436 N_A_1175_93#_c_655_n N_A_1004_379#_M1007_g 0.00203946f $X=7.08 $Y=1.615
+ $X2=0 $Y2=0
cc_437 N_A_1175_93#_M1001_g N_A_1004_379#_c_740_n 0.00214917f $X=5.95 $Y=0.805
+ $X2=0 $Y2=0
cc_438 N_A_1175_93#_M1001_g N_A_1004_379#_c_741_n 0.0117608f $X=5.95 $Y=0.805
+ $X2=0 $Y2=0
cc_439 N_A_1175_93#_c_644_n N_A_1004_379#_c_741_n 0.0191306f $X=6.1 $Y=1.725
+ $X2=0 $Y2=0
cc_440 N_A_1175_93#_c_652_n N_A_1004_379#_c_741_n 0.00979f $X=6.75 $Y=1.72 $X2=0
+ $Y2=0
cc_441 N_A_1175_93#_c_664_n N_A_1004_379#_c_741_n 0.0236023f $X=6.19 $Y=1.56
+ $X2=0 $Y2=0
cc_442 N_A_1175_93#_c_644_n N_A_1004_379#_c_742_n 0.00555599f $X=6.1 $Y=1.725
+ $X2=0 $Y2=0
cc_443 N_A_1175_93#_c_664_n N_A_1004_379#_c_742_n 0.013704f $X=6.19 $Y=1.56
+ $X2=0 $Y2=0
cc_444 N_A_1175_93#_c_644_n N_A_1004_379#_c_743_n 0.00120939f $X=6.1 $Y=1.725
+ $X2=0 $Y2=0
cc_445 N_A_1175_93#_c_652_n N_A_1004_379#_c_743_n 0.0127092f $X=6.75 $Y=1.72
+ $X2=0 $Y2=0
cc_446 N_A_1175_93#_c_653_n N_A_1004_379#_c_743_n 0.0221035f $X=7.08 $Y=1.425
+ $X2=0 $Y2=0
cc_447 N_A_1175_93#_c_654_n N_A_1004_379#_c_743_n 0.0078729f $X=6.855 $Y=0.52
+ $X2=0 $Y2=0
cc_448 N_A_1175_93#_c_655_n N_A_1004_379#_c_743_n 0.00840588f $X=7.08 $Y=1.615
+ $X2=0 $Y2=0
cc_449 N_A_1175_93#_c_644_n N_A_1004_379#_c_744_n 0.0312278f $X=6.1 $Y=1.725
+ $X2=0 $Y2=0
cc_450 N_A_1175_93#_c_649_n N_A_1004_379#_c_744_n 0.00684647f $X=7.63 $Y=1.51
+ $X2=0 $Y2=0
cc_451 N_A_1175_93#_c_652_n N_A_1004_379#_c_744_n 2.41424e-19 $X=6.75 $Y=1.72
+ $X2=0 $Y2=0
cc_452 N_A_1175_93#_c_653_n N_A_1004_379#_c_744_n 0.00584137f $X=7.08 $Y=1.425
+ $X2=0 $Y2=0
cc_453 N_A_1175_93#_c_654_n N_A_1004_379#_c_744_n 0.00367342f $X=6.855 $Y=0.52
+ $X2=0 $Y2=0
cc_454 N_A_1175_93#_c_655_n N_A_1004_379#_c_744_n 0.00390355f $X=7.08 $Y=1.615
+ $X2=0 $Y2=0
cc_455 N_A_1175_93#_M1001_g N_A_1004_379#_c_745_n 0.00903736f $X=5.95 $Y=0.805
+ $X2=0 $Y2=0
cc_456 N_A_1175_93#_c_653_n N_A_1004_379#_c_745_n 0.00439627f $X=7.08 $Y=1.425
+ $X2=0 $Y2=0
cc_457 N_A_1175_93#_c_654_n N_A_1004_379#_c_745_n 0.00617551f $X=6.855 $Y=0.52
+ $X2=0 $Y2=0
cc_458 N_A_1175_93#_c_644_n N_VPWR_c_819_n 9.98489e-19 $X=6.1 $Y=1.725 $X2=0
+ $Y2=0
cc_459 N_A_1175_93#_M1020_g N_VPWR_c_819_n 0.0106716f $X=6.1 $Y=2.105 $X2=0
+ $Y2=0
cc_460 N_A_1175_93#_c_652_n N_VPWR_c_819_n 0.0134455f $X=6.75 $Y=1.72 $X2=0
+ $Y2=0
cc_461 N_A_1175_93#_c_663_n N_VPWR_c_819_n 0.00135677f $X=6.855 $Y=2.04 $X2=0
+ $Y2=0
cc_462 N_A_1175_93#_c_664_n N_VPWR_c_819_n 0.0149433f $X=6.19 $Y=1.56 $X2=0
+ $Y2=0
cc_463 N_A_1175_93#_M1008_g N_VPWR_c_820_n 0.00767118f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_464 N_A_1175_93#_c_649_n N_VPWR_c_820_n 0.00776673f $X=7.63 $Y=1.51 $X2=0
+ $Y2=0
cc_465 N_A_1175_93#_c_663_n N_VPWR_c_820_n 0.0786911f $X=6.855 $Y=2.04 $X2=0
+ $Y2=0
cc_466 N_A_1175_93#_c_655_n N_VPWR_c_820_n 0.00816477f $X=7.08 $Y=1.615 $X2=0
+ $Y2=0
cc_467 N_A_1175_93#_M1019_g N_VPWR_c_822_n 0.00770354f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_A_1175_93#_c_663_n N_VPWR_c_827_n 0.00952375f $X=6.855 $Y=2.04 $X2=0
+ $Y2=0
cc_469 N_A_1175_93#_M1008_g N_VPWR_c_828_n 0.00585385f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_470 N_A_1175_93#_M1019_g N_VPWR_c_828_n 0.00585385f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_471 N_A_1175_93#_M1020_g N_VPWR_c_814_n 0.00314105f $X=6.1 $Y=2.105 $X2=0
+ $Y2=0
cc_472 N_A_1175_93#_M1008_g N_VPWR_c_814_n 0.0118358f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_473 N_A_1175_93#_M1019_g N_VPWR_c_814_n 0.0114822f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_474 N_A_1175_93#_c_663_n N_VPWR_c_814_n 0.0130956f $X=6.855 $Y=2.04 $X2=0
+ $Y2=0
cc_475 N_A_1175_93#_c_645_n Q 0.00239621f $X=7.705 $Y=1.345 $X2=0 $Y2=0
cc_476 N_A_1175_93#_c_646_n Q 0.018333f $X=8.06 $Y=1.42 $X2=0 $Y2=0
cc_477 N_A_1175_93#_c_647_n Q 0.00352479f $X=8.135 $Y=1.345 $X2=0 $Y2=0
cc_478 N_A_1175_93#_M1019_g Q 0.00948635f $X=8.135 $Y=2.465 $X2=0 $Y2=0
cc_479 N_A_1175_93#_c_650_n Q 0.00522617f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_480 N_A_1175_93#_c_663_n Q 3.17794e-19 $X=6.855 $Y=2.04 $X2=0 $Y2=0
cc_481 N_A_1175_93#_c_653_n Q 0.00472603f $X=7.08 $Y=1.425 $X2=0 $Y2=0
cc_482 N_A_1175_93#_c_655_n Q 0.0154017f $X=7.08 $Y=1.615 $X2=0 $Y2=0
cc_483 N_A_1175_93#_M1001_g N_VGND_c_964_n 0.0112638f $X=5.95 $Y=0.805 $X2=0
+ $Y2=0
cc_484 N_A_1175_93#_c_644_n N_VGND_c_964_n 0.00178928f $X=6.1 $Y=1.725 $X2=0
+ $Y2=0
cc_485 N_A_1175_93#_c_645_n N_VGND_c_965_n 0.00742594f $X=7.705 $Y=1.345 $X2=0
+ $Y2=0
cc_486 N_A_1175_93#_c_649_n N_VGND_c_965_n 0.00828997f $X=7.63 $Y=1.51 $X2=0
+ $Y2=0
cc_487 N_A_1175_93#_c_654_n N_VGND_c_965_n 0.0690625f $X=6.855 $Y=0.52 $X2=0
+ $Y2=0
cc_488 N_A_1175_93#_c_655_n N_VGND_c_965_n 0.00816421f $X=7.08 $Y=1.615 $X2=0
+ $Y2=0
cc_489 N_A_1175_93#_c_647_n N_VGND_c_967_n 0.00742395f $X=8.135 $Y=1.345 $X2=0
+ $Y2=0
cc_490 N_A_1175_93#_M1001_g N_VGND_c_971_n 0.0035863f $X=5.95 $Y=0.805 $X2=0
+ $Y2=0
cc_491 N_A_1175_93#_c_654_n N_VGND_c_972_n 0.0152962f $X=6.855 $Y=0.52 $X2=0
+ $Y2=0
cc_492 N_A_1175_93#_c_645_n N_VGND_c_973_n 0.00559701f $X=7.705 $Y=1.345 $X2=0
+ $Y2=0
cc_493 N_A_1175_93#_c_647_n N_VGND_c_973_n 0.00559701f $X=8.135 $Y=1.345 $X2=0
+ $Y2=0
cc_494 N_A_1175_93#_M1001_g N_VGND_c_976_n 0.00401353f $X=5.95 $Y=0.805 $X2=0
+ $Y2=0
cc_495 N_A_1175_93#_c_645_n N_VGND_c_976_n 0.00537853f $X=7.705 $Y=1.345 $X2=0
+ $Y2=0
cc_496 N_A_1175_93#_c_647_n N_VGND_c_976_n 0.00537853f $X=8.135 $Y=1.345 $X2=0
+ $Y2=0
cc_497 N_A_1175_93#_c_654_n N_VGND_c_976_n 0.0165373f $X=6.855 $Y=0.52 $X2=0
+ $Y2=0
cc_498 N_A_1004_379#_M1007_g N_VPWR_c_819_n 0.00773706f $X=6.64 $Y=2.315 $X2=0
+ $Y2=0
cc_499 N_A_1004_379#_c_748_n N_VPWR_c_819_n 0.0224942f $X=5.43 $Y=2.04 $X2=0
+ $Y2=0
cc_500 N_A_1004_379#_M1007_g N_VPWR_c_820_n 0.0035373f $X=6.64 $Y=2.315 $X2=0
+ $Y2=0
cc_501 N_A_1004_379#_c_748_n N_VPWR_c_823_n 0.00733305f $X=5.43 $Y=2.04 $X2=0
+ $Y2=0
cc_502 N_A_1004_379#_M1007_g N_VPWR_c_827_n 0.00431487f $X=6.64 $Y=2.315 $X2=0
+ $Y2=0
cc_503 N_A_1004_379#_M1007_g N_VPWR_c_814_n 0.00477801f $X=6.64 $Y=2.315 $X2=0
+ $Y2=0
cc_504 N_A_1004_379#_c_748_n N_VPWR_c_814_n 0.0100833f $X=5.43 $Y=2.04 $X2=0
+ $Y2=0
cc_505 N_A_1004_379#_c_740_n N_VGND_c_964_n 0.013698f $X=5.57 $Y=1.295 $X2=0
+ $Y2=0
cc_506 N_A_1004_379#_c_741_n N_VGND_c_964_n 0.03796f $X=6.565 $Y=1.21 $X2=0
+ $Y2=0
cc_507 N_A_1004_379#_c_745_n N_VGND_c_964_n 0.00768951f $X=6.73 $Y=1.125 $X2=0
+ $Y2=0
cc_508 N_A_1004_379#_c_745_n N_VGND_c_965_n 0.00345282f $X=6.73 $Y=1.125 $X2=0
+ $Y2=0
cc_509 N_A_1004_379#_c_740_n N_VGND_c_971_n 0.00869096f $X=5.57 $Y=1.295 $X2=0
+ $Y2=0
cc_510 N_A_1004_379#_c_745_n N_VGND_c_972_n 0.00431792f $X=6.73 $Y=1.125 $X2=0
+ $Y2=0
cc_511 N_A_1004_379#_c_740_n N_VGND_c_976_n 0.0130067f $X=5.57 $Y=1.295 $X2=0
+ $Y2=0
cc_512 N_A_1004_379#_c_745_n N_VGND_c_976_n 0.00544287f $X=6.73 $Y=1.125 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_814_n N_Q_M1008_d 0.0027574f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_514 N_VPWR_c_820_n Q 0.00153572f $X=7.49 $Y=1.98 $X2=0 $Y2=0
cc_515 N_VPWR_c_822_n Q 0.00151552f $X=8.35 $Y=1.98 $X2=0 $Y2=0
cc_516 N_VPWR_c_828_n Q 0.0151136f $X=8.22 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_c_814_n Q 0.0102248f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_518 N_VPWR_c_820_n N_VGND_c_965_n 0.00720482f $X=7.49 $Y=1.98 $X2=0 $Y2=0
cc_519 N_VPWR_c_822_n N_VGND_c_967_n 0.0094937f $X=8.35 $Y=1.98 $X2=0 $Y2=0
cc_520 N_A_432_119#_c_919_n N_VGND_c_963_n 0.0235228f $X=2.53 $Y=0.805 $X2=0
+ $Y2=0
cc_521 N_A_432_119#_c_919_n N_VGND_c_970_n 0.00663586f $X=2.53 $Y=0.805 $X2=0
+ $Y2=0
cc_522 N_A_432_119#_c_919_n N_VGND_c_976_n 0.00996178f $X=2.53 $Y=0.805 $X2=0
+ $Y2=0
cc_523 Q N_VGND_c_965_n 0.00307144f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_524 Q N_VGND_c_967_n 0.00303104f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_525 Q N_VGND_c_973_n 0.0106634f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_526 Q N_VGND_c_976_n 0.00956577f $X=7.835 $Y=0.47 $X2=0 $Y2=0
