* File: sky130_fd_sc_lp__o211a_1.pxi.spice
* Created: Wed Sep  2 10:13:45 2020
* 
x_PM_SKY130_FD_SC_LP__O211A_1%A_80_237# N_A_80_237#_M1009_d N_A_80_237#_M1001_d
+ N_A_80_237#_M1006_d N_A_80_237#_c_59_n N_A_80_237#_M1003_g N_A_80_237#_M1007_g
+ N_A_80_237#_c_111_p N_A_80_237#_c_61_n N_A_80_237#_c_62_n N_A_80_237#_c_63_n
+ N_A_80_237#_c_75_p N_A_80_237#_c_119_p N_A_80_237#_c_125_p N_A_80_237#_c_93_p
+ N_A_80_237#_c_64_n N_A_80_237#_c_68_n N_A_80_237#_c_69_n N_A_80_237#_c_65_n
+ N_A_80_237#_c_89_p PM_SKY130_FD_SC_LP__O211A_1%A_80_237#
x_PM_SKY130_FD_SC_LP__O211A_1%A1 N_A1_M1004_g N_A1_M1000_g A1 N_A1_c_153_n
+ N_A1_c_156_n PM_SKY130_FD_SC_LP__O211A_1%A1
x_PM_SKY130_FD_SC_LP__O211A_1%A2 N_A2_M1001_g N_A2_M1005_g A2 N_A2_c_190_n
+ N_A2_c_193_n PM_SKY130_FD_SC_LP__O211A_1%A2
x_PM_SKY130_FD_SC_LP__O211A_1%B1 N_B1_M1002_g N_B1_M1008_g B1 B1 N_B1_c_225_n
+ PM_SKY130_FD_SC_LP__O211A_1%B1
x_PM_SKY130_FD_SC_LP__O211A_1%C1 N_C1_M1009_g N_C1_M1006_g N_C1_c_258_n C1
+ N_C1_c_259_n N_C1_c_260_n PM_SKY130_FD_SC_LP__O211A_1%C1
x_PM_SKY130_FD_SC_LP__O211A_1%X N_X_M1003_s N_X_M1007_s X X X X X X X
+ N_X_c_284_n X N_X_c_287_n PM_SKY130_FD_SC_LP__O211A_1%X
x_PM_SKY130_FD_SC_LP__O211A_1%VPWR N_VPWR_M1007_d N_VPWR_M1002_d N_VPWR_c_303_n
+ N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n VPWR N_VPWR_c_307_n
+ N_VPWR_c_308_n N_VPWR_c_302_n N_VPWR_c_310_n PM_SKY130_FD_SC_LP__O211A_1%VPWR
x_PM_SKY130_FD_SC_LP__O211A_1%VGND N_VGND_M1003_d N_VGND_M1004_d N_VGND_c_345_n
+ N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n VGND N_VGND_c_349_n
+ N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n PM_SKY130_FD_SC_LP__O211A_1%VGND
x_PM_SKY130_FD_SC_LP__O211A_1%A_266_49# N_A_266_49#_M1004_s N_A_266_49#_M1005_d
+ N_A_266_49#_c_392_n N_A_266_49#_c_397_n N_A_266_49#_c_393_n
+ N_A_266_49#_c_401_n N_A_266_49#_c_419_n PM_SKY130_FD_SC_LP__O211A_1%A_266_49#
cc_1 VNB N_A_80_237#_c_59_n 0.0222277f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.185
cc_2 VNB N_A_80_237#_M1007_g 0.00930611f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_3 VNB N_A_80_237#_c_61_n 0.0747798f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.35
cc_4 VNB N_A_80_237#_c_62_n 0.00234937f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.92
cc_5 VNB N_A_80_237#_c_63_n 0.0351044f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.11
cc_6 VNB N_A_80_237#_c_64_n 0.0300527f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=0.42
cc_7 VNB N_A_80_237#_c_65_n 0.014934f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.27
cc_8 VNB N_A1_M1004_g 0.031129f $X=-0.19 $Y=-0.245 $X2=3.265 $Y2=1.835
cc_9 VNB N_A1_c_153_n 0.0279088f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.655
cc_10 VNB N_A2_M1005_g 0.0274906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_190_n 0.0257481f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.655
cc_12 VNB N_B1_M1008_g 0.0238865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB B1 0.00410321f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.185
cc_14 VNB N_B1_c_225_n 0.0220411f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_15 VNB N_C1_M1009_g 0.0268061f $X=-0.19 $Y=-0.245 $X2=3.265 $Y2=1.835
cc_16 VNB N_C1_M1006_g 0.00138783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C1_c_258_n 0.00909218f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.185
cc_18 VNB N_C1_c_259_n 0.0540061f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_19 VNB N_C1_c_260_n 0.0126243f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_20 VNB X 0.0406294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_284_n 0.0247063f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.11
cc_22 VNB N_VPWR_c_302_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_345_n 0.0133673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_346_n 0.00602232f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.52
cc_25 VNB N_VGND_c_347_n 0.0245699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_348_n 0.00631736f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.35
cc_27 VNB N_VGND_c_349_n 0.0166266f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.35
cc_28 VNB N_VGND_c_350_n 0.0487684f $X=-0.19 $Y=-0.245 $X2=2.545 $Y2=2.005
cc_29 VNB N_VGND_c_351_n 0.231961f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=1.025
cc_30 VNB N_VGND_c_352_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_266_49#_c_392_n 0.00539916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_266_49#_c_393_n 0.00242156f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.655
cc_33 VPB N_A_80_237#_M1007_g 0.0272982f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.465
cc_34 VPB N_A_80_237#_c_62_n 0.00446299f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.92
cc_35 VPB N_A_80_237#_c_68_n 0.00743679f $X=-0.19 $Y=1.655 $X2=3.41 $Y2=2.09
cc_36 VPB N_A_80_237#_c_69_n 0.0382376f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=2.91
cc_37 VPB N_A1_M1000_g 0.0205787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A1_c_153_n 0.00663762f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.655
cc_39 VPB N_A1_c_156_n 0.00219186f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.52
cc_40 VPB N_A2_M1001_g 0.0192409f $X=-0.19 $Y=1.655 $X2=3.265 $Y2=1.835
cc_41 VPB N_A2_c_190_n 0.00647396f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.655
cc_42 VPB N_A2_c_193_n 0.00211949f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.52
cc_43 VPB N_B1_M1002_g 0.0208218f $X=-0.19 $Y=1.655 $X2=3.265 $Y2=1.835
cc_44 VPB B1 0.00462894f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.185
cc_45 VPB N_B1_c_225_n 0.00613159f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.465
cc_46 VPB N_C1_M1006_g 0.0262782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_C1_c_260_n 0.0128605f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.465
cc_48 VPB X 0.00940833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB X 0.0574151f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.655
cc_50 VPB N_X_c_287_n 0.0309563f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.352
cc_51 VPB N_VPWR_c_303_n 0.00192478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_304_n 0.0055721f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.52
cc_53 VPB N_VPWR_c_305_n 0.029217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_306_n 0.00631825f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.35
cc_55 VPB N_VPWR_c_307_n 0.026601f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.35
cc_56 VPB N_VPWR_c_308_n 0.0232155f $X=-0.19 $Y=1.655 $X2=2.38 $Y2=2.475
cc_57 VPB N_VPWR_c_302_n 0.056054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_310_n 0.0104351f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=1.025
cc_59 N_A_80_237#_c_61_n N_A1_M1004_g 0.00280701f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_60 N_A_80_237#_c_63_n N_A1_M1004_g 0.0130734f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_61 N_A_80_237#_c_65_n N_A1_M1004_g 0.00394812f $X=1.205 $Y=1.27 $X2=0 $Y2=0
cc_62 N_A_80_237#_M1007_g N_A1_M1000_g 0.0107034f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A_80_237#_c_62_n N_A1_M1000_g 0.00362923f $X=1.205 $Y=1.92 $X2=0 $Y2=0
cc_64 N_A_80_237#_c_75_p N_A1_M1000_g 0.0149947f $X=2.215 $Y=2.005 $X2=0 $Y2=0
cc_65 N_A_80_237#_M1007_g N_A1_c_153_n 0.00296224f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_80_237#_c_61_n N_A1_c_153_n 0.00447662f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_67 N_A_80_237#_c_62_n N_A1_c_153_n 0.00132236f $X=1.205 $Y=1.92 $X2=0 $Y2=0
cc_68 N_A_80_237#_c_63_n N_A1_c_153_n 0.00448227f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_69 N_A_80_237#_c_75_p N_A1_c_153_n 9.19902e-19 $X=2.215 $Y=2.005 $X2=0 $Y2=0
cc_70 N_A_80_237#_c_65_n N_A1_c_153_n 0.00188067f $X=1.205 $Y=1.27 $X2=0 $Y2=0
cc_71 N_A_80_237#_c_62_n N_A1_c_156_n 0.018407f $X=1.205 $Y=1.92 $X2=0 $Y2=0
cc_72 N_A_80_237#_c_63_n N_A1_c_156_n 0.0245052f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_73 N_A_80_237#_c_75_p N_A1_c_156_n 0.022946f $X=2.215 $Y=2.005 $X2=0 $Y2=0
cc_74 N_A_80_237#_c_65_n N_A1_c_156_n 0.01265f $X=1.205 $Y=1.27 $X2=0 $Y2=0
cc_75 N_A_80_237#_c_75_p N_A2_M1001_g 0.0124277f $X=2.215 $Y=2.005 $X2=0 $Y2=0
cc_76 N_A_80_237#_c_63_n N_A2_M1005_g 0.0118338f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_77 N_A_80_237#_c_63_n N_A2_c_190_n 0.00474865f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_78 N_A_80_237#_c_89_p N_A2_c_190_n 8.88922e-19 $X=2.38 $Y=2.005 $X2=0 $Y2=0
cc_79 N_A_80_237#_c_63_n N_A2_c_193_n 0.024509f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_80 N_A_80_237#_c_75_p N_A2_c_193_n 0.0120804f $X=2.215 $Y=2.005 $X2=0 $Y2=0
cc_81 N_A_80_237#_c_89_p N_A2_c_193_n 0.011908f $X=2.38 $Y=2.005 $X2=0 $Y2=0
cc_82 N_A_80_237#_c_93_p N_B1_M1002_g 0.0135135f $X=3.25 $Y=2.005 $X2=0 $Y2=0
cc_83 N_A_80_237#_c_69_n N_B1_M1002_g 7.29221e-19 $X=3.405 $Y=2.91 $X2=0 $Y2=0
cc_84 N_A_80_237#_c_63_n N_B1_M1008_g 0.0150921f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_85 N_A_80_237#_c_64_n N_B1_M1008_g 0.00253269f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_86 N_A_80_237#_c_63_n B1 0.0511099f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_87 N_A_80_237#_c_93_p B1 0.0452425f $X=3.25 $Y=2.005 $X2=0 $Y2=0
cc_88 N_A_80_237#_c_63_n N_B1_c_225_n 0.00473543f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_89 N_A_80_237#_c_93_p N_B1_c_225_n 9.21682e-19 $X=3.25 $Y=2.005 $X2=0 $Y2=0
cc_90 N_A_80_237#_c_63_n N_C1_M1009_g 0.0155813f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_91 N_A_80_237#_c_64_n N_C1_M1009_g 0.015853f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_80_237#_c_93_p N_C1_M1006_g 0.0137513f $X=3.25 $Y=2.005 $X2=0 $Y2=0
cc_93 N_A_80_237#_c_68_n N_C1_M1006_g 9.50925e-19 $X=3.41 $Y=2.09 $X2=0 $Y2=0
cc_94 N_A_80_237#_c_69_n N_C1_M1006_g 0.0136896f $X=3.405 $Y=2.91 $X2=0 $Y2=0
cc_95 N_A_80_237#_c_63_n N_C1_c_259_n 0.0104437f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_96 N_A_80_237#_c_68_n N_C1_c_259_n 0.00455148f $X=3.41 $Y=2.09 $X2=0 $Y2=0
cc_97 N_A_80_237#_c_63_n N_C1_c_260_n 0.0157571f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_98 N_A_80_237#_c_68_n N_C1_c_260_n 0.0162788f $X=3.41 $Y=2.09 $X2=0 $Y2=0
cc_99 N_A_80_237#_c_59_n X 0.00611857f $X=0.535 $Y=1.185 $X2=0 $Y2=0
cc_100 N_A_80_237#_c_111_p X 0.0269166f $X=1.085 $Y=1.35 $X2=0 $Y2=0
cc_101 N_A_80_237#_c_61_n X 0.0171723f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_102 N_A_80_237#_M1007_g N_X_c_287_n 0.00338927f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_80_237#_c_111_p N_X_c_287_n 0.0198426f $X=1.085 $Y=1.35 $X2=0 $Y2=0
cc_104 N_A_80_237#_c_61_n N_X_c_287_n 0.0121421f $X=0.925 $Y=1.35 $X2=0 $Y2=0
cc_105 N_A_80_237#_c_62_n N_X_c_287_n 0.00134349f $X=1.205 $Y=1.92 $X2=0 $Y2=0
cc_106 N_A_80_237#_c_62_n N_VPWR_M1007_d 0.00215484f $X=1.205 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_80_237#_c_75_p N_VPWR_M1007_d 0.0122094f $X=2.215 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_108 N_A_80_237#_c_119_p N_VPWR_M1007_d 0.00428275f $X=1.325 $Y=2.005
+ $X2=-0.19 $Y2=-0.245
cc_109 N_A_80_237#_c_93_p N_VPWR_M1002_d 0.00590163f $X=3.25 $Y=2.005 $X2=0
+ $Y2=0
cc_110 N_A_80_237#_M1007_g N_VPWR_c_303_n 0.0201724f $X=0.98 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_80_237#_c_75_p N_VPWR_c_303_n 0.0255877f $X=2.215 $Y=2.005 $X2=0
+ $Y2=0
cc_112 N_A_80_237#_c_119_p N_VPWR_c_303_n 0.0191594f $X=1.325 $Y=2.005 $X2=0
+ $Y2=0
cc_113 N_A_80_237#_c_93_p N_VPWR_c_304_n 0.022455f $X=3.25 $Y=2.005 $X2=0 $Y2=0
cc_114 N_A_80_237#_c_125_p N_VPWR_c_305_n 0.0212513f $X=2.38 $Y=2.475 $X2=0
+ $Y2=0
cc_115 N_A_80_237#_M1007_g N_VPWR_c_307_n 0.00486043f $X=0.98 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_80_237#_c_69_n N_VPWR_c_308_n 0.0203649f $X=3.405 $Y=2.91 $X2=0 $Y2=0
cc_117 N_A_80_237#_M1001_d N_VPWR_c_302_n 0.00521751f $X=2.185 $Y=1.835 $X2=0
+ $Y2=0
cc_118 N_A_80_237#_M1006_d N_VPWR_c_302_n 0.00215158f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_119 N_A_80_237#_M1007_g N_VPWR_c_302_n 0.00954696f $X=0.98 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_80_237#_c_125_p N_VPWR_c_302_n 0.0127519f $X=2.38 $Y=2.475 $X2=0
+ $Y2=0
cc_121 N_A_80_237#_c_69_n N_VPWR_c_302_n 0.0122259f $X=3.405 $Y=2.91 $X2=0 $Y2=0
cc_122 N_A_80_237#_c_75_p A_365_367# 0.00732587f $X=2.215 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_80_237#_c_63_n N_VGND_M1004_d 0.0041528f $X=3.24 $Y=1.11 $X2=0 $Y2=0
cc_124 N_A_80_237#_c_59_n N_VGND_c_345_n 0.0181975f $X=0.535 $Y=1.185 $X2=0
+ $Y2=0
cc_125 N_A_80_237#_c_111_p N_VGND_c_345_n 0.0244884f $X=1.085 $Y=1.35 $X2=0
+ $Y2=0
cc_126 N_A_80_237#_c_61_n N_VGND_c_345_n 0.00694369f $X=0.925 $Y=1.35 $X2=0
+ $Y2=0
cc_127 N_A_80_237#_c_59_n N_VGND_c_349_n 0.00486043f $X=0.535 $Y=1.185 $X2=0
+ $Y2=0
cc_128 N_A_80_237#_c_64_n N_VGND_c_350_n 0.0210467f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_129 N_A_80_237#_M1009_d N_VGND_c_351_n 0.00212301f $X=3.265 $Y=0.245 $X2=0
+ $Y2=0
cc_130 N_A_80_237#_c_59_n N_VGND_c_351_n 0.00923188f $X=0.535 $Y=1.185 $X2=0
+ $Y2=0
cc_131 N_A_80_237#_c_64_n N_VGND_c_351_n 0.0125689f $X=3.405 $Y=0.42 $X2=0 $Y2=0
cc_132 N_A_80_237#_c_63_n N_A_266_49#_M1004_s 0.00248866f $X=3.24 $Y=1.11
+ $X2=-0.19 $Y2=-0.245
cc_133 N_A_80_237#_c_63_n N_A_266_49#_M1005_d 0.0030319f $X=3.24 $Y=1.11 $X2=0
+ $Y2=0
cc_134 N_A_80_237#_c_59_n N_A_266_49#_c_392_n 0.00111122f $X=0.535 $Y=1.185
+ $X2=0 $Y2=0
cc_135 N_A_80_237#_c_63_n N_A_266_49#_c_397_n 0.0444293f $X=3.24 $Y=1.11 $X2=0
+ $Y2=0
cc_136 N_A_80_237#_c_59_n N_A_266_49#_c_393_n 5.22876e-19 $X=0.535 $Y=1.185
+ $X2=0 $Y2=0
cc_137 N_A_80_237#_c_63_n N_A_266_49#_c_393_n 0.018975f $X=3.24 $Y=1.11 $X2=0
+ $Y2=0
cc_138 N_A_80_237#_c_65_n N_A_266_49#_c_393_n 0.00324972f $X=1.205 $Y=1.27 $X2=0
+ $Y2=0
cc_139 N_A_80_237#_c_63_n N_A_266_49#_c_401_n 0.0222271f $X=3.24 $Y=1.11 $X2=0
+ $Y2=0
cc_140 N_A_80_237#_c_63_n A_581_49# 0.00366293f $X=3.24 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A1_M1000_g N_A2_M1001_g 0.0569745f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A1_M1004_g N_A2_M1005_g 0.0290725f $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_143 N_A1_c_153_n N_A2_c_190_n 0.0569745f $X=1.66 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A1_c_156_n N_A2_c_190_n 0.00130275f $X=1.66 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A1_c_153_n N_A2_c_193_n 0.00130275f $X=1.66 $Y=1.51 $X2=0 $Y2=0
cc_146 N_A1_c_156_n N_A2_c_193_n 0.0243354f $X=1.66 $Y=1.51 $X2=0 $Y2=0
cc_147 N_A1_M1000_g N_VPWR_c_303_n 0.0240733f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A1_M1000_g N_VPWR_c_305_n 0.00486043f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A1_M1000_g N_VPWR_c_302_n 0.00818711f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A1_M1004_g N_VGND_c_345_n 0.0040274f $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_151 N_A1_M1004_g N_VGND_c_346_n 0.00585742f $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_152 N_A1_M1004_g N_VGND_c_347_n 0.00413177f $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_153 N_A1_M1004_g N_VGND_c_351_n 0.00753387f $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_154 N_A1_M1004_g N_A_266_49#_c_392_n 0.00661421f $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_155 N_A1_M1004_g N_A_266_49#_c_397_n 0.00950756f $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_156 N_A1_M1004_g N_A_266_49#_c_393_n 7.15802e-19 $X=1.67 $Y=0.665 $X2=0 $Y2=0
cc_157 N_A2_M1001_g N_B1_M1002_g 0.0133234f $X=2.11 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A2_c_193_n N_B1_M1002_g 2.55411e-19 $X=2.2 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A2_M1005_g N_B1_M1008_g 0.0172552f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_160 N_A2_M1001_g B1 2.0934e-19 $X=2.11 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A2_c_190_n B1 0.00187963f $X=2.2 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A2_c_193_n B1 0.0325641f $X=2.2 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A2_c_190_n N_B1_c_225_n 0.0208742f $X=2.2 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A2_c_193_n N_B1_c_225_n 3.55575e-19 $X=2.2 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A2_M1001_g N_VPWR_c_303_n 0.00357156f $X=2.11 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A2_M1001_g N_VPWR_c_305_n 0.00585385f $X=2.11 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A2_M1001_g N_VPWR_c_302_n 0.0109726f $X=2.11 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_M1005_g N_VGND_c_346_n 0.00608829f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_169 N_A2_M1005_g N_VGND_c_350_n 0.00423815f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_170 N_A2_M1005_g N_VGND_c_351_n 0.00662677f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_171 N_A2_M1005_g N_A_266_49#_c_392_n 8.05532e-19 $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_172 N_A2_M1005_g N_A_266_49#_c_397_n 0.0108503f $X=2.29 $Y=0.665 $X2=0 $Y2=0
cc_173 N_B1_M1008_g N_C1_M1009_g 0.0486124f $X=2.83 $Y=0.665 $X2=0 $Y2=0
cc_174 N_B1_M1002_g N_C1_M1006_g 0.0324426f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_175 B1 N_C1_M1006_g 0.00471854f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_176 B1 N_C1_c_258_n 0.00970704f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_177 N_B1_c_225_n N_C1_c_258_n 0.0486124f $X=2.74 $Y=1.51 $X2=0 $Y2=0
cc_178 B1 N_C1_c_260_n 0.0298829f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B1_M1002_g N_VPWR_c_304_n 0.00441125f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B1_M1002_g N_VPWR_c_305_n 0.00585385f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B1_M1002_g N_VPWR_c_302_n 0.0110984f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B1_M1008_g N_VGND_c_350_n 0.00575161f $X=2.83 $Y=0.665 $X2=0 $Y2=0
cc_183 N_B1_M1008_g N_VGND_c_351_n 0.0109364f $X=2.83 $Y=0.665 $X2=0 $Y2=0
cc_184 N_C1_M1006_g N_VPWR_c_304_n 0.00804767f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_185 N_C1_M1006_g N_VPWR_c_308_n 0.00564131f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_186 N_C1_M1006_g N_VPWR_c_302_n 0.0115657f $X=3.19 $Y=2.465 $X2=0 $Y2=0
cc_187 N_C1_M1009_g N_VGND_c_350_n 0.00539298f $X=3.19 $Y=0.665 $X2=0 $Y2=0
cc_188 N_C1_M1009_g N_VGND_c_351_n 0.0108778f $X=3.19 $Y=0.665 $X2=0 $Y2=0
cc_189 X N_VPWR_c_307_n 0.0547298f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_190 N_X_M1007_s N_VPWR_c_302_n 0.00371702f $X=0.64 $Y=1.835 $X2=0 $Y2=0
cc_191 X N_VPWR_c_302_n 0.0300525f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_192 X N_VGND_c_345_n 8.05345e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_193 N_X_c_284_n N_VGND_c_349_n 0.0228292f $X=0.32 $Y=0.42 $X2=0 $Y2=0
cc_194 N_X_M1003_s N_VGND_c_351_n 0.00371702f $X=0.195 $Y=0.235 $X2=0 $Y2=0
cc_195 N_X_c_284_n N_VGND_c_351_n 0.0127519f $X=0.32 $Y=0.42 $X2=0 $Y2=0
cc_196 N_VPWR_c_302_n A_365_367# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_197 N_VGND_c_351_n N_A_266_49#_M1004_s 0.00212301f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_198 N_VGND_c_351_n N_A_266_49#_M1005_d 0.00428094f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_345_n N_A_266_49#_c_392_n 0.020702f $X=0.75 $Y=0.38 $X2=0 $Y2=0
cc_200 N_VGND_c_346_n N_A_266_49#_c_392_n 0.0181582f $X=1.98 $Y=0.41 $X2=0 $Y2=0
cc_201 N_VGND_c_347_n N_A_266_49#_c_392_n 0.0208729f $X=1.815 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_351_n N_A_266_49#_c_392_n 0.0125275f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_M1004_d N_A_266_49#_c_397_n 0.00847899f $X=1.745 $Y=0.245 $X2=0
+ $Y2=0
cc_204 N_VGND_c_346_n N_A_266_49#_c_397_n 0.0253821f $X=1.98 $Y=0.41 $X2=0 $Y2=0
cc_205 N_VGND_c_347_n N_A_266_49#_c_397_n 0.00250142f $X=1.815 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_350_n N_A_266_49#_c_397_n 0.00312364f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_351_n N_A_266_49#_c_397_n 0.0122187f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_208 N_VGND_c_345_n N_A_266_49#_c_393_n 0.00868461f $X=0.75 $Y=0.38 $X2=0
+ $Y2=0
cc_209 N_VGND_c_350_n N_A_266_49#_c_419_n 0.0210745f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_351_n N_A_266_49#_c_419_n 0.0127102f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_351_n A_581_49# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
