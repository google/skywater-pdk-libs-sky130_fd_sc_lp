* NGSPICE file created from sky130_fd_sc_lp__dlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
M1000 a_1078_367# CLK VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=2.7749e+12p ps=1.959e+07u
M1001 a_73_269# a_295_55# a_253_81# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1002 a_1078_367# a_27_367# a_1026_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=1.764e+11p ps=2.1e+06u
M1003 VPWR a_1078_367# GCLK VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1004 GCLK a_1078_367# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=1.46918e+12p ps=1.352e+07u
M1005 a_1026_47# CLK VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_235_465# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1007 a_415_465# a_295_55# a_73_269# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.221e+11p ps=2.06e+06u
M1008 a_277_367# a_295_55# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 a_253_81# GATE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_27_367# a_411_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1011 VPWR a_27_367# a_415_465# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR CLK a_295_55# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.7485e+11p ps=2.21e+06u
M1013 VGND a_1078_367# GCLK VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_411_81# a_277_367# a_73_269# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_1078_367# GCLK VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 GCLK a_1078_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_27_367# a_1078_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 GCLK a_1078_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 GCLK a_1078_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_73_269# a_277_367# a_235_465# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_277_367# a_295_55# VPWR VPB phighvt w=640000u l=150000u
+  ad=2.25e+11p pd=2.03e+06u as=0p ps=0u
M1022 VGND a_73_269# a_27_367# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1023 VPWR a_1078_367# GCLK VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND CLK a_295_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.999e+11p ps=1.86e+06u
M1025 VPWR a_73_269# a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

