* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buf_m A VGND VNB VPB VPWR X
X0 X a_47_178# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_47_178# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND A a_47_178# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR A a_47_178# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
