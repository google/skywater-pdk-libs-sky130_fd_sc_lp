* File: sky130_fd_sc_lp__o311a_4.pex.spice
* Created: Fri Aug 28 11:13:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311A_4%A_81_23# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 54 57 61 63 65 66 69 73 75 77 81 94
c129 75 0 1.7348e-19 $X=5.122 $Y=1.875
r130 91 92 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.715 $Y=1.49
+ $X2=1.77 $Y2=1.49
r131 90 91 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.34 $Y=1.49
+ $X2=1.715 $Y2=1.49
r132 89 90 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.285 $Y=1.49
+ $X2=1.34 $Y2=1.49
r133 88 89 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.91 $Y=1.49
+ $X2=1.285 $Y2=1.49
r134 87 88 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.855 $Y=1.49
+ $X2=0.91 $Y2=1.49
r135 75 83 3.0159 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=5.122 $Y=1.875
+ $X2=5.122 $Y2=1.79
r136 75 77 35.5977 $w=2.23e-07 $l=6.95e-07 $layer=LI1_cond $X=5.122 $Y=1.875
+ $X2=5.122 $Y2=2.57
r137 74 81 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.82 $Y=1.79
+ $X2=3.707 $Y2=1.79
r138 73 83 3.9739 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=5.01 $Y=1.79
+ $X2=5.122 $Y2=1.79
r139 73 74 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=5.01 $Y=1.79
+ $X2=3.82 $Y2=1.79
r140 69 71 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=3.707 $Y=1.98
+ $X2=3.707 $Y2=2.91
r141 67 81 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.707 $Y=1.875
+ $X2=3.707 $Y2=1.79
r142 67 69 5.37807 $w=2.23e-07 $l=1.05e-07 $layer=LI1_cond $X=3.707 $Y=1.875
+ $X2=3.707 $Y2=1.98
r143 65 81 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.595 $Y=1.79
+ $X2=3.707 $Y2=1.79
r144 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.595 $Y=1.79
+ $X2=2.925 $Y2=1.79
r145 61 63 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=2.795 $Y=0.89
+ $X2=2.935 $Y2=0.89
r146 57 59 46.5988 $w=2.28e-07 $l=9.3e-07 $layer=LI1_cond $X=2.81 $Y=1.98
+ $X2=2.81 $Y2=2.91
r147 55 66 7.76265 $w=4.16e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.81 $Y=1.875
+ $X2=2.925 $Y2=1.79
r148 55 57 5.26115 $w=2.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.81 $Y=1.875
+ $X2=2.81 $Y2=1.98
r149 54 55 7.41971 $w=4.16e-07 $l=3.51374e-07 $layer=LI1_cond $X=2.557 $Y=1.64
+ $X2=2.81 $Y2=1.875
r150 53 61 7.70722 $w=2.5e-07 $l=2.93929e-07 $layer=LI1_cond $X=2.557 $Y=1.015
+ $X2=2.795 $Y2=0.89
r151 53 54 9.82043 $w=4.73e-07 $l=3.9e-07 $layer=LI1_cond $X=2.557 $Y=1.015
+ $X2=2.557 $Y2=1.405
r152 52 94 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.055 $Y=1.49
+ $X2=2.145 $Y2=1.49
r153 52 92 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.055 $Y=1.49
+ $X2=1.77 $Y2=1.49
r154 51 52 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.055
+ $Y=1.49 $X2=2.055 $Y2=1.49
r155 48 87 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.695 $Y=1.49
+ $X2=0.855 $Y2=1.49
r156 48 84 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.695 $Y=1.49
+ $X2=0.48 $Y2=1.49
r157 47 51 83.798 $w=1.78e-07 $l=1.36e-06 $layer=LI1_cond $X=0.695 $Y=1.495
+ $X2=2.055 $Y2=1.495
r158 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.695
+ $Y=1.49 $X2=0.695 $Y2=1.49
r159 45 54 14.6168 $w=4.16e-07 $l=4.28409e-07 $layer=LI1_cond $X=2.195 $Y=1.495
+ $X2=2.557 $Y2=1.64
r160 45 51 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.195 $Y=1.495
+ $X2=2.055 $Y2=1.495
r161 41 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.655
+ $X2=2.145 $Y2=1.49
r162 41 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.145 $Y=1.655
+ $X2=2.145 $Y2=2.465
r163 37 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=1.49
r164 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.77 $Y=1.325
+ $X2=1.77 $Y2=0.665
r165 33 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.655
+ $X2=1.715 $Y2=1.49
r166 33 35 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.715 $Y=1.655
+ $X2=1.715 $Y2=2.465
r167 29 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=1.49
r168 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.34 $Y=1.325
+ $X2=1.34 $Y2=0.665
r169 25 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.655
+ $X2=1.285 $Y2=1.49
r170 25 27 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.285 $Y=1.655
+ $X2=1.285 $Y2=2.465
r171 21 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.49
r172 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=0.665
r173 17 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.855 $Y=1.655
+ $X2=0.855 $Y2=1.49
r174 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.855 $Y=1.655
+ $X2=0.855 $Y2=2.465
r175 13 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.49
r176 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=0.665
r177 4 83 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.725 $X2=5.105 $Y2=1.87
r178 4 77 400 $w=1.7e-07 $l=9.12318e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.725 $X2=5.105 $Y2=2.57
r179 3 71 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.835 $X2=3.725 $Y2=2.91
r180 3 69 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.835 $X2=3.725 $Y2=1.98
r181 2 59 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.835 $X2=2.79 $Y2=2.91
r182 2 57 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.835 $X2=2.79 $Y2=1.98
r183 1 63 182 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.235 $X2=2.935 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%C1 3 5 7 10 12 14 15 21
r46 21 23 14.3642 $w=3.02e-07 $l=9e-08 $layer=POLY_cond $X=3.06 $Y=1.355
+ $X2=3.15 $Y2=1.355
r47 19 21 8.77815 $w=3.02e-07 $l=5.5e-08 $layer=POLY_cond $X=3.005 $Y=1.355
+ $X2=3.06 $Y2=1.355
r48 18 19 45.4868 $w=3.02e-07 $l=2.85e-07 $layer=POLY_cond $X=2.72 $Y=1.355
+ $X2=3.005 $Y2=1.355
r49 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.36 $X2=3.06 $Y2=1.36
r50 12 23 19.1248 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.15 $Y=1.185
+ $X2=3.15 $Y2=1.355
r51 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.15 $Y=1.185
+ $X2=3.15 $Y2=0.655
r52 8 19 19.1248 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.005 $Y=1.525
+ $X2=3.005 $Y2=1.355
r53 8 10 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.005 $Y=1.525 $X2=3.005
+ $Y2=2.465
r54 5 18 19.1248 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.72 $Y=1.185
+ $X2=2.72 $Y2=1.355
r55 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.72 $Y=1.185 $X2=2.72
+ $Y2=0.655
r56 1 18 23.1424 $w=3.02e-07 $l=2.31409e-07 $layer=POLY_cond $X=2.575 $Y=1.525
+ $X2=2.72 $Y2=1.355
r57 1 3 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.575 $Y=1.525 $X2=2.575
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%B1 3 5 7 10 12 14 15 24
c43 24 0 1.46531e-19 $X=4.01 $Y=1.385
r44 23 24 10.2449 $w=3.8e-07 $l=7e-08 $layer=POLY_cond $X=3.94 $Y=1.385 $X2=4.01
+ $Y2=1.385
r45 21 23 49.7611 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=3.6 $Y=1.385
+ $X2=3.94 $Y2=1.385
r46 19 21 2.92713 $w=3.8e-07 $l=2e-08 $layer=POLY_cond $X=3.58 $Y=1.385 $X2=3.6
+ $Y2=1.385
r47 17 19 10.2449 $w=3.8e-07 $l=7e-08 $layer=POLY_cond $X=3.51 $Y=1.385 $X2=3.58
+ $Y2=1.385
r48 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=1.36 $X2=3.6 $Y2=1.36
r49 12 24 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.01 $Y=1.195
+ $X2=4.01 $Y2=1.385
r50 12 14 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.01 $Y=1.195
+ $X2=4.01 $Y2=0.655
r51 8 23 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.94 $Y=1.575
+ $X2=3.94 $Y2=1.385
r52 8 10 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.94 $Y=1.575
+ $X2=3.94 $Y2=2.465
r53 5 19 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.58 $Y=1.195
+ $X2=3.58 $Y2=1.385
r54 5 7 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.58 $Y=1.195 $X2=3.58
+ $Y2=0.655
r55 1 17 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.51 $Y=1.575
+ $X2=3.51 $Y2=1.385
r56 1 3 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.51 $Y=1.575 $X2=3.51
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%A3 3 5 7 10 12 14 15 20 21 22 23 24
c51 24 0 4.23065e-20 $X=5.52 $Y=1.295
c52 20 0 1.13451e-19 $X=5.815 $Y=1.35
c53 10 0 1.7348e-19 $X=5.32 $Y=2.355
r54 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.41
+ $Y=1.35 $X2=5.41 $Y2=1.35
r55 24 31 4.15635 $w=3.03e-07 $l=1.1e-07 $layer=LI1_cond $X=5.52 $Y=1.362
+ $X2=5.41 $Y2=1.362
r56 23 31 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=5.04 $Y=1.362
+ $X2=5.41 $Y2=1.362
r57 22 23 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.362
+ $X2=5.04 $Y2=1.362
r58 21 22 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.362
+ $X2=4.56 $Y2=1.362
r59 20 30 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=5.815 $Y=1.35
+ $X2=5.41 $Y2=1.35
r60 18 19 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.96 $Y=1.35
+ $X2=5.32 $Y2=1.35
r61 16 18 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.89 $Y=1.35 $X2=4.96
+ $Y2=1.35
r62 15 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.395 $Y=1.35
+ $X2=5.41 $Y2=1.35
r63 15 19 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.395 $Y=1.35
+ $X2=5.32 $Y2=1.35
r64 12 20 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.89 $Y=1.185
+ $X2=5.815 $Y2=1.35
r65 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.89 $Y=1.185
+ $X2=5.89 $Y2=0.655
r66 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.515
+ $X2=5.32 $Y2=1.35
r67 8 10 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.32 $Y=1.515
+ $X2=5.32 $Y2=2.355
r68 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.96 $Y=1.185
+ $X2=4.96 $Y2=1.35
r69 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.96 $Y=1.185 $X2=4.96
+ $Y2=0.655
r70 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.515
+ $X2=4.89 $Y2=1.35
r71 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.89 $Y=1.515 $X2=4.89
+ $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%A2 3 7 11 15 17 18 19 28
c56 28 0 1.96579e-19 $X=6.75 $Y=1.51
c57 19 0 5.82438e-20 $X=6.96 $Y=1.665
r58 26 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.41 $Y=1.51
+ $X2=6.75 $Y2=1.51
r59 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=1.51 $X2=6.41 $Y2=1.51
r60 23 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.32 $Y=1.51 $X2=6.41
+ $Y2=1.51
r61 18 19 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.592
+ $X2=6.96 $Y2=1.592
r62 18 27 2.40809 $w=3.33e-07 $l=7e-08 $layer=LI1_cond $X=6.48 $Y=1.592 $X2=6.41
+ $Y2=1.592
r63 17 27 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=6 $Y=1.592 $X2=6.41
+ $Y2=1.592
r64 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.75 $Y=1.675
+ $X2=6.75 $Y2=1.51
r65 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.75 $Y=1.675
+ $X2=6.75 $Y2=2.465
r66 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.75 $Y=1.345
+ $X2=6.75 $Y2=1.51
r67 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.75 $Y=1.345
+ $X2=6.75 $Y2=0.655
r68 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.32 $Y=1.675
+ $X2=6.32 $Y2=1.51
r69 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.32 $Y=1.675 $X2=6.32
+ $Y2=2.465
r70 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.32 $Y=1.345
+ $X2=6.32 $Y2=1.51
r71 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.32 $Y=1.345 $X2=6.32
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%A1 3 7 11 15 17 18 26
c38 18 0 1.54272e-19 $X=7.92 $Y=1.665
c39 15 0 5.82438e-20 $X=7.61 $Y=2.465
r40 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.52 $Y=1.51 $X2=7.61
+ $Y2=1.51
r41 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.52
+ $Y=1.51 $X2=7.52 $Y2=1.51
r42 21 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.18 $Y=1.51
+ $X2=7.52 $Y2=1.51
r43 18 25 13.7605 $w=3.33e-07 $l=4e-07 $layer=LI1_cond $X=7.92 $Y=1.592 $X2=7.52
+ $Y2=1.592
r44 17 25 2.7521 $w=3.33e-07 $l=8e-08 $layer=LI1_cond $X=7.44 $Y=1.592 $X2=7.52
+ $Y2=1.592
r45 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.61 $Y=1.675
+ $X2=7.61 $Y2=1.51
r46 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.61 $Y=1.675
+ $X2=7.61 $Y2=2.465
r47 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.61 $Y=1.345
+ $X2=7.61 $Y2=1.51
r48 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.61 $Y=1.345
+ $X2=7.61 $Y2=0.655
r49 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.18 $Y=1.675
+ $X2=7.18 $Y2=1.51
r50 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.18 $Y=1.675 $X2=7.18
+ $Y2=2.465
r51 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.18 $Y=1.345
+ $X2=7.18 $Y2=1.51
r52 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.18 $Y=1.345 $X2=7.18
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%VPWR 1 2 3 4 5 6 21 27 33 37 41 47 53 56 57
+ 58 59 60 62 74 79 89 90 93 96 99 102
r109 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r111 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 90 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 87 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.56 $Y=3.33
+ $X2=7.395 $Y2=3.33
r115 87 89 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.56 $Y=3.33
+ $X2=7.92 $Y2=3.33
r116 86 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r117 85 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 83 86 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 82 85 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.96 $Y2=3.33
r120 82 83 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r121 80 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.155 $Y2=3.33
r122 80 82 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r123 79 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=3.33
+ $X2=7.395 $Y2=3.33
r124 79 85 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.23 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r127 75 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r128 75 77 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 74 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=4.155 $Y2=3.33
r130 74 77 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=3.6 $Y2=3.33
r131 73 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r133 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r134 70 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r135 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r136 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.64 $Y2=3.33
r137 67 69 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 65 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 62 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.64 $Y2=3.33
r141 62 64 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.24 $Y2=3.33
r142 60 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 60 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r144 60 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 58 72 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.16 $Y2=3.33
r146 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.36 $Y2=3.33
r147 56 69 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.5 $Y2=3.33
r149 55 72 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=2.16 $Y2=3.33
r150 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=1.5 $Y2=3.33
r151 51 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=3.245
+ $X2=7.395 $Y2=3.33
r152 51 53 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=7.395 $Y=3.245
+ $X2=7.395 $Y2=2.39
r153 47 50 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.155 $Y=2.13
+ $X2=4.155 $Y2=2.95
r154 45 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=3.33
r155 45 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=2.95
r156 41 44 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=3.26 $Y=2.13
+ $X2=3.26 $Y2=2.95
r157 39 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r158 39 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.95
r159 38 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.36 $Y2=3.33
r160 37 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r161 37 38 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=2.525 $Y2=3.33
r162 33 36 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=2.36 $Y=2.13
+ $X2=2.36 $Y2=2.95
r163 31 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=3.245
+ $X2=2.36 $Y2=3.33
r164 31 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=3.245
+ $X2=2.36 $Y2=2.95
r165 27 30 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.5 $Y=2.19 $X2=1.5
+ $Y2=2.95
r166 25 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=3.245 $X2=1.5
+ $Y2=3.33
r167 25 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.5 $Y=3.245
+ $X2=1.5 $Y2=2.95
r168 21 24 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.64 $Y=2.18
+ $X2=0.64 $Y2=2.95
r169 19 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=3.245
+ $X2=0.64 $Y2=3.33
r170 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.64 $Y=3.245
+ $X2=0.64 $Y2=2.95
r171 6 53 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=7.255
+ $Y=1.835 $X2=7.395 $Y2=2.39
r172 5 50 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.835 $X2=4.155 $Y2=2.95
r173 5 47 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.835 $X2=4.155 $Y2=2.13
r174 4 44 400 $w=1.7e-07 $l=1.20163e-06 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.835 $X2=3.26 $Y2=2.95
r175 4 41 400 $w=1.7e-07 $l=3.74333e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.835 $X2=3.26 $Y2=2.13
r176 3 36 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.835 $X2=2.36 $Y2=2.95
r177 3 33 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=1.835 $X2=2.36 $Y2=2.13
r178 2 30 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.95
r179 2 27 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.19
r180 1 24 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.515
+ $Y=1.835 $X2=0.64 $Y2=2.95
r181 1 21 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.515
+ $Y=1.835 $X2=0.64 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%X 1 2 3 4 13 15 16 19 21 25 29 33 37 42 43
+ 44 45 49 51
r56 49 51 2.51442 $w=2.73e-07 $l=6e-08 $layer=LI1_cond $X=0.222 $Y=1.235
+ $X2=0.222 $Y2=1.295
r57 44 49 2.84615 $w=2.75e-07 $l=9e-08 $layer=LI1_cond $X=0.222 $Y=1.145
+ $X2=0.222 $Y2=1.235
r58 44 45 15.0027 $w=2.73e-07 $l=3.58e-07 $layer=LI1_cond $X=0.222 $Y=1.307
+ $X2=0.222 $Y2=1.665
r59 44 51 0.502884 $w=2.73e-07 $l=1.2e-08 $layer=LI1_cond $X=0.222 $Y=1.307
+ $X2=0.222 $Y2=1.295
r60 41 45 3.77163 $w=2.73e-07 $l=9e-08 $layer=LI1_cond $X=0.222 $Y=1.755
+ $X2=0.222 $Y2=1.665
r61 37 39 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.93 $Y=1.98
+ $X2=1.93 $Y2=2.91
r62 35 37 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.93 $Y=1.925
+ $X2=1.93 $Y2=1.98
r63 31 33 32.3185 $w=2.28e-07 $l=6.45e-07 $layer=LI1_cond $X=1.575 $Y=1.065
+ $X2=1.575 $Y2=0.42
r64 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.165 $Y=1.84
+ $X2=1.07 $Y2=1.84
r65 29 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.835 $Y=1.84
+ $X2=1.93 $Y2=1.925
r66 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.835 $Y=1.84
+ $X2=1.165 $Y2=1.84
r67 25 27 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.07 $Y=1.98
+ $X2=1.07 $Y2=2.91
r68 23 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=1.925
+ $X2=1.07 $Y2=1.84
r69 23 25 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.07 $Y=1.925
+ $X2=1.07 $Y2=1.98
r70 22 42 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=0.79 $Y=1.15
+ $X2=0.695 $Y2=1.145
r71 21 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.46 $Y=1.15
+ $X2=1.575 $Y2=1.065
r72 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.46 $Y=1.15
+ $X2=0.79 $Y2=1.15
r73 17 42 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=0.695 $Y=1.055
+ $X2=0.695 $Y2=1.145
r74 17 19 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.695 $Y=1.055
+ $X2=0.695 $Y2=0.42
r75 16 41 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=0.36 $Y=1.84
+ $X2=0.222 $Y2=1.755
r76 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.975 $Y=1.84
+ $X2=1.07 $Y2=1.84
r77 15 16 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.975 $Y=1.84
+ $X2=0.36 $Y2=1.84
r78 14 44 4.3641 $w=1.8e-07 $l=1.38e-07 $layer=LI1_cond $X=0.36 $Y=1.145
+ $X2=0.222 $Y2=1.145
r79 13 42 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=0.6 $Y=1.145
+ $X2=0.695 $Y2=1.145
r80 13 14 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.6 $Y=1.145
+ $X2=0.36 $Y2=1.145
r81 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=2.91
r82 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.835 $X2=1.93 $Y2=1.98
r83 3 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=1.835 $X2=1.07 $Y2=2.91
r84 3 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=1.835 $X2=1.07 $Y2=1.98
r85 2 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.415
+ $Y=0.245 $X2=1.555 $Y2=0.42
r86 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.245 $X2=0.695 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%A_910_345# 1 2 3 12 16 17 20 24 28 30
r43 26 28 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.535 $Y=2.905
+ $X2=6.535 $Y2=2.39
r44 25 30 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.68 $Y=2.99
+ $X2=5.542 $Y2=2.99
r45 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.37 $Y=2.99
+ $X2=6.535 $Y2=2.905
r46 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.37 $Y=2.99 $X2=5.68
+ $Y2=2.99
r47 20 23 40.6498 $w=2.73e-07 $l=9.7e-07 $layer=LI1_cond $X=5.542 $Y=1.87
+ $X2=5.542 $Y2=2.84
r48 18 30 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.542 $Y=2.905
+ $X2=5.542 $Y2=2.99
r49 18 23 2.72396 $w=2.73e-07 $l=6.5e-08 $layer=LI1_cond $X=5.542 $Y=2.905
+ $X2=5.542 $Y2=2.84
r50 16 30 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=5.405 $Y=2.99
+ $X2=5.542 $Y2=2.99
r51 16 17 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.405 $Y=2.99
+ $X2=4.84 $Y2=2.99
r52 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.675 $Y=2.13
+ $X2=4.675 $Y2=2.84
r53 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.675 $Y=2.905
+ $X2=4.84 $Y2=2.99
r54 10 15 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=4.675 $Y=2.905
+ $X2=4.675 $Y2=2.84
r55 3 28 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=6.395
+ $Y=1.835 $X2=6.535 $Y2=2.39
r56 2 23 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.725 $X2=5.535 $Y2=2.84
r57 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.725 $X2=5.535 $Y2=1.87
r58 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=4.55
+ $Y=1.725 $X2=4.675 $Y2=2.84
r59 1 12 400 $w=1.7e-07 $l=4.63303e-07 $layer=licon1_PDIFF $count=1 $X=4.55
+ $Y=1.725 $X2=4.675 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%A_1196_367# 1 2 3 10 12 14 18 20 22 24 29
c32 10 0 1.13451e-19 $X=6.07 $Y=2.1
r33 22 31 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=2.1 $X2=7.86
+ $Y2=2.015
r34 22 24 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=7.86 $Y=2.1 $X2=7.86
+ $Y2=2.45
r35 21 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.06 $Y=2.015
+ $X2=6.965 $Y2=2.015
r36 20 31 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.73 $Y=2.015
+ $X2=7.86 $Y2=2.015
r37 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.73 $Y=2.015
+ $X2=7.06 $Y2=2.015
r38 16 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=2.1
+ $X2=6.965 $Y2=2.015
r39 16 18 19.555 $w=1.88e-07 $l=3.35e-07 $layer=LI1_cond $X=6.965 $Y=2.1
+ $X2=6.965 $Y2=2.435
r40 15 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.2 $Y=2.015 $X2=6.07
+ $Y2=2.015
r41 14 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.87 $Y=2.015
+ $X2=6.965 $Y2=2.015
r42 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.87 $Y=2.015
+ $X2=6.2 $Y2=2.015
r43 10 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=2.1 $X2=6.07
+ $Y2=2.015
r44 10 12 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=6.07 $Y=2.1 $X2=6.07
+ $Y2=2.57
r45 3 31 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.835 $X2=7.825 $Y2=2.015
r46 3 24 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=7.685
+ $Y=1.835 $X2=7.825 $Y2=2.45
r47 2 29 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=6.825
+ $Y=1.835 $X2=6.965 $Y2=2.015
r48 2 18 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=6.825
+ $Y=1.835 $X2=6.965 $Y2=2.435
r49 1 27 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=5.98
+ $Y=1.835 $X2=6.105 $Y2=2.015
r50 1 12 600 $w=1.7e-07 $l=7.95047e-07 $layer=licon1_PDIFF $count=1 $X=5.98
+ $Y=1.835 $X2=6.105 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 40 41 42
+ 44 57 62 69 70 76 81 87 89 92
r112 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r113 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r114 86 87 11.3415 $w=7.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=0.307
+ $X2=5.84 $Y2=0.307
r115 83 86 2.36168 $w=7.83e-07 $l=1.55e-07 $layer=LI1_cond $X=5.52 $Y=0.307
+ $X2=5.675 $Y2=0.307
r116 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r117 80 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r118 79 83 7.3136 $w=7.83e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=0.307
+ $X2=5.52 $Y2=0.307
r119 79 81 9.28454 $w=7.83e-07 $l=3e-08 $layer=LI1_cond $X=5.04 $Y=0.307
+ $X2=5.01 $Y2=0.307
r120 79 80 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r121 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r122 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 70 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r124 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r125 67 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.56 $Y=0 $X2=7.395
+ $Y2=0
r126 67 69 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.56 $Y=0 $X2=7.92
+ $Y2=0
r127 66 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r128 66 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r129 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r130 63 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.7 $Y=0 $X2=6.535
+ $Y2=0
r131 63 65 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.7 $Y=0 $X2=6.96
+ $Y2=0
r132 62 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=0 $X2=7.395
+ $Y2=0
r133 62 65 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.23 $Y=0 $X2=6.96
+ $Y2=0
r134 61 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r135 61 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r136 60 87 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6 $Y=0 $X2=5.84
+ $Y2=0
r137 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r138 57 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6.535
+ $Y2=0
r139 57 60 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6
+ $Y2=0
r140 55 81 185.936 $w=1.68e-07 $l=2.85e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=5.01
+ $Y2=0
r141 55 56 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r142 52 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r143 52 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r144 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r145 49 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.125
+ $Y2=0
r146 49 51 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.68
+ $Y2=0
r147 48 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r148 48 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r149 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r150 45 73 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r151 45 47 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r152 44 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.125
+ $Y2=0
r153 44 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r154 42 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r155 42 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.16 $Y2=0
r156 40 51 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.68
+ $Y2=0
r157 40 41 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.005
+ $Y2=0
r158 39 55 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.16
+ $Y2=0
r159 39 41 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.005
+ $Y2=0
r160 35 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=0.085
+ $X2=7.395 $Y2=0
r161 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.395 $Y=0.085
+ $X2=7.395 $Y2=0.38
r162 31 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=0.085
+ $X2=6.535 $Y2=0
r163 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.535 $Y=0.085
+ $X2=6.535 $Y2=0.38
r164 27 41 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0
r165 27 29 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0.39
r166 23 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0
r167 23 25 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.125 $Y=0.085
+ $X2=1.125 $Y2=0.37
r168 19 73 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.215 $Y2=0
r169 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.39
r170 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.255
+ $Y=0.235 $X2=7.395 $Y2=0.38
r171 5 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.395
+ $Y=0.235 $X2=6.535 $Y2=0.38
r172 4 86 91 $w=1.7e-07 $l=7.87909e-07 $layer=licon1_NDIFF $count=2 $X=5.035
+ $Y=0.235 $X2=5.675 $Y2=0.565
r173 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.845
+ $Y=0.245 $X2=1.985 $Y2=0.39
r174 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.245 $X2=1.125 $Y2=0.37
r175 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.245 $X2=0.265 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%A_476_47# 1 2 3 10 16 18 21 22
c31 16 0 1.46531e-19 $X=3.365 $Y=0.86
r32 22 25 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=4.26 $Y=0.345
+ $X2=4.26 $Y2=0.52
r33 19 21 3.9502 $w=2.6e-07 $l=1.28938e-07 $layer=LI1_cond $X=3.46 $Y=0.345
+ $X2=3.365 $Y2=0.425
r34 18 22 2.89065 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.13 $Y=0.345
+ $X2=4.26 $Y2=0.345
r35 18 19 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.13 $Y=0.345
+ $X2=3.46 $Y2=0.345
r36 14 21 2.49283 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=3.365 $Y=0.595
+ $X2=3.365 $Y2=0.425
r37 14 16 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=3.365 $Y=0.595
+ $X2=3.365 $Y2=0.86
r38 10 21 3.9502 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=3.27 $Y=0.425
+ $X2=3.365 $Y2=0.425
r39 10 12 25.93 $w=3.38e-07 $l=7.65e-07 $layer=LI1_cond $X=3.27 $Y=0.425
+ $X2=2.505 $Y2=0.425
r40 3 25 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=4.085
+ $Y=0.235 $X2=4.225 $Y2=0.52
r41 2 21 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.235 $X2=3.365 $Y2=0.42
r42 2 16 182 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.235 $X2=3.365 $Y2=0.86
r43 1 12 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.505 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O311A_4%A_731_47# 1 2 3 4 5 16 20 22 26 28 32 34 38
+ 41 43 44 48
c66 32 0 1.37393e-19 $X=6.965 $Y=0.42
r67 44 46 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=6.1 $Y=0.955
+ $X2=6.1 $Y2=1.17
r68 44 45 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=6.1 $Y=0.955 $X2=6.1
+ $Y2=0.87
r69 41 42 7.17421 $w=3.18e-07 $l=1.87e-07 $layer=LI1_cond $X=3.795 $Y=0.76
+ $X2=3.795 $Y2=0.947
r70 36 38 29.4759 $w=2.58e-07 $l=6.65e-07 $layer=LI1_cond $X=7.86 $Y=1.085
+ $X2=7.86 $Y2=0.42
r71 35 48 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.06 $Y=1.17
+ $X2=6.965 $Y2=1.17
r72 34 36 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.73 $Y=1.17
+ $X2=7.86 $Y2=1.085
r73 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.73 $Y=1.17
+ $X2=7.06 $Y2=1.17
r74 30 48 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=1.085
+ $X2=6.965 $Y2=1.17
r75 30 32 38.8182 $w=1.88e-07 $l=6.65e-07 $layer=LI1_cond $X=6.965 $Y=1.085
+ $X2=6.965 $Y2=0.42
r76 29 46 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.2 $Y=1.17 $X2=6.1
+ $Y2=1.17
r77 28 48 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.87 $Y=1.17
+ $X2=6.965 $Y2=1.17
r78 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.87 $Y=1.17 $X2=6.2
+ $Y2=1.17
r79 26 45 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=6.105 $Y=0.42
+ $X2=6.105 $Y2=0.87
r80 23 43 7.00709 $w=1.77e-07 $l=1.3394e-07 $layer=LI1_cond $X=4.84 $Y=0.955
+ $X2=4.71 $Y2=0.947
r81 22 44 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6 $Y=0.955 $X2=6.1
+ $Y2=0.955
r82 22 23 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=6 $Y=0.955 $X2=4.84
+ $Y2=0.955
r83 18 43 0.0115521 $w=2.6e-07 $l=9.2e-08 $layer=LI1_cond $X=4.71 $Y=0.855
+ $X2=4.71 $Y2=0.947
r84 18 20 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=4.71 $Y=0.855
+ $X2=4.71 $Y2=0.42
r85 17 42 3.92581 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=3.96 $Y=0.947
+ $X2=3.795 $Y2=0.947
r86 16 43 7.00709 $w=1.77e-07 $l=1.3e-07 $layer=LI1_cond $X=4.58 $Y=0.947
+ $X2=4.71 $Y2=0.947
r87 16 17 37.1695 $w=1.83e-07 $l=6.2e-07 $layer=LI1_cond $X=4.58 $Y=0.947
+ $X2=3.96 $Y2=0.947
r88 5 38 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.685
+ $Y=0.235 $X2=7.825 $Y2=0.42
r89 4 32 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.825
+ $Y=0.235 $X2=6.965 $Y2=0.42
r90 3 26 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.965
+ $Y=0.235 $X2=6.105 $Y2=0.42
r91 2 20 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=4.62
+ $Y=0.235 $X2=4.745 $Y2=0.42
r92 1 41 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.235 $X2=3.795 $Y2=0.76
.ends

