# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__xor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.260000 1.180000 1.550000 1.225000 ;
        RECT 1.260000 1.225000 6.625000 1.365000 ;
        RECT 1.260000 1.365000 1.550000 1.410000 ;
        RECT 3.455000 1.180000 3.745000 1.225000 ;
        RECT 3.455000 1.365000 3.745000 1.410000 ;
        RECT 6.335000 1.180000 6.625000 1.225000 ;
        RECT 6.335000 1.365000 6.625000 1.410000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.495000 1.550000 2.785000 1.595000 ;
        RECT 2.495000 1.595000 8.065000 1.735000 ;
        RECT 2.495000 1.735000 2.785000 1.780000 ;
        RECT 7.775000 1.550000 8.065000 1.595000 ;
        RECT 7.775000 1.735000 8.065000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815000 0.695000 4.295000 0.905000 ;
        RECT 3.995000 0.905000 4.295000 1.015000 ;
        RECT 3.995000 1.015000 5.155000 1.185000 ;
        RECT 3.995000 1.185000 4.275000 2.290000 ;
        RECT 3.995000 2.290000 5.195000 2.605000 ;
        RECT 4.105000 0.255000 4.295000 0.695000 ;
        RECT 4.865000 1.845000 5.195000 2.290000 ;
        RECT 4.965000 0.255000 5.155000 1.015000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.095000  0.085000  0.425000 1.095000 ;
      RECT 0.095000  1.695000  1.225000 1.865000 ;
      RECT 0.095000  1.865000  0.355000 3.075000 ;
      RECT 0.400000  1.275000  1.555000 1.525000 ;
      RECT 0.525000  2.035000  0.855000 3.245000 ;
      RECT 0.595000  0.255000  0.815000 0.735000 ;
      RECT 0.595000  0.735000  1.645000 0.905000 ;
      RECT 0.595000  0.905000  0.785000 1.095000 ;
      RECT 0.985000  0.085000  1.215000 0.565000 ;
      RECT 1.025000  1.865000  1.225000 1.945000 ;
      RECT 1.025000  1.945000  3.825000 2.115000 ;
      RECT 1.025000  2.115000  1.215000 3.075000 ;
      RECT 1.260000  1.075000  3.685000 1.245000 ;
      RECT 1.260000  1.245000  1.555000 1.275000 ;
      RECT 1.385000  0.255000  3.435000 0.525000 ;
      RECT 1.385000  0.525000  1.645000 0.735000 ;
      RECT 1.385000  2.285000  1.715000 3.245000 ;
      RECT 1.735000  1.415000  3.085000 1.775000 ;
      RECT 1.885000  2.115000  2.075000 3.075000 ;
      RECT 2.245000  2.285000  2.575000 3.245000 ;
      RECT 2.745000  2.115000  2.950000 3.075000 ;
      RECT 3.120000  2.285000  3.450000 3.245000 ;
      RECT 3.340000  1.245000  3.685000 1.435000 ;
      RECT 3.605000  0.085000  3.935000 0.525000 ;
      RECT 3.625000  2.115000  3.825000 2.775000 ;
      RECT 3.625000  2.775000  5.625000 3.075000 ;
      RECT 4.445000  1.355000  6.135000 1.535000 ;
      RECT 4.465000  0.085000  4.795000 0.845000 ;
      RECT 5.325000  0.085000  6.215000 0.690000 ;
      RECT 5.325000  0.690000  5.655000 1.105000 ;
      RECT 5.365000  1.815000  5.625000 2.775000 ;
      RECT 5.825000  0.860000  7.435000 1.015000 ;
      RECT 5.825000  1.015000  9.995000 1.030000 ;
      RECT 5.825000  1.030000  6.135000 1.355000 ;
      RECT 5.955000  1.970000  7.935000 2.140000 ;
      RECT 5.955000  2.140000  6.215000 3.075000 ;
      RECT 6.305000  1.200000  7.075000 1.355000 ;
      RECT 6.305000  1.355000  7.655000 1.535000 ;
      RECT 6.385000  0.255000  6.575000 0.860000 ;
      RECT 6.385000  2.310000  6.715000 3.245000 ;
      RECT 6.745000  0.085000  7.075000 0.690000 ;
      RECT 6.885000  2.140000  7.075000 3.075000 ;
      RECT 7.245000  0.255000  7.435000 0.860000 ;
      RECT 7.245000  1.030000  9.995000 1.185000 ;
      RECT 7.245000  2.310000  7.575000 3.245000 ;
      RECT 7.605000  0.085000  7.935000 0.845000 ;
      RECT 7.745000  2.140000  7.935000 2.905000 ;
      RECT 7.745000  2.905000  9.725000 3.075000 ;
      RECT 7.825000  1.355000  9.600000 1.535000 ;
      RECT 7.825000  1.535000  8.015000 1.800000 ;
      RECT 8.105000  0.255000  8.295000 1.015000 ;
      RECT 8.185000  1.705000  9.995000 1.875000 ;
      RECT 8.185000  1.875000  8.435000 2.735000 ;
      RECT 8.465000  0.085000  8.795000 0.845000 ;
      RECT 8.605000  2.045000  8.795000 2.905000 ;
      RECT 8.965000  0.255000  9.155000 1.015000 ;
      RECT 8.965000  1.875000  9.295000 2.735000 ;
      RECT 9.325000  0.085000  9.655000 0.845000 ;
      RECT 9.465000  2.045000  9.725000 2.905000 ;
      RECT 9.770000  1.185000  9.995000 1.705000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.320000  1.210000 1.490000 1.380000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.580000 2.725000 1.750000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  1.210000 3.685000 1.380000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  1.210000 6.565000 1.380000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  1.580000 8.005000 1.750000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__xor2_4
END LIBRARY
