* File: sky130_fd_sc_lp__sdfrtp_ov2.pex.spice
* Created: Fri Aug 28 11:28:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_35_74# 1 2 7 9 12 15 18 21 22 24 26 31
+ 33 34 41
c73 33 0 8.22072e-20 $X=2.51 $Y=1.98
c74 22 0 1.42315e-19 $X=1.345 $Y=0.945
r75 34 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.98
+ $X2=2.51 $Y2=2.145
r76 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.98 $X2=2.51 $Y2=1.98
r77 30 31 12.3626 $w=9.88e-07 $l=1.3e-07 $layer=LI1_cond $X=1.01 $Y=2.47
+ $X2=1.14 $Y2=2.47
r78 27 30 9.61212 $w=9.88e-07 $l=7.8e-07 $layer=LI1_cond $X=0.23 $Y=2.47
+ $X2=1.01 $Y2=2.47
r79 24 33 2.99516 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=2.425 $Y=2.06
+ $X2=2.55 $Y2=1.98
r80 24 31 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=2.425 $Y=2.06
+ $X2=1.14 $Y2=2.06
r81 22 38 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=1.345 $Y=0.945
+ $X2=1.465 $Y2=0.945
r82 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=0.945 $X2=1.345 $Y2=0.945
r83 19 26 3.57226 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.43 $Y=0.945
+ $X2=0.26 $Y2=0.945
r84 19 21 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=0.43 $Y=0.945
+ $X2=1.345 $Y2=0.945
r85 18 27 8.32829 $w=2.8e-07 $l=4.95e-07 $layer=LI1_cond $X=0.23 $Y=1.975
+ $X2=0.23 $Y2=2.47
r86 17 26 3.05675 $w=3.1e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.23 $Y=1.03
+ $X2=0.26 $Y2=0.945
r87 17 18 38.895 $w=2.78e-07 $l=9.45e-07 $layer=LI1_cond $X=0.23 $Y=1.03
+ $X2=0.23 $Y2=1.975
r88 13 26 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.86 $X2=0.26
+ $Y2=0.945
r89 13 15 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=0.26 $Y=0.86
+ $X2=0.26 $Y2=0.58
r90 12 41 122.107 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.49 $Y=2.525
+ $X2=2.49 $Y2=2.145
r91 7 38 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=0.78
+ $X2=1.465 $Y2=0.945
r92 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.465 $Y=0.78
+ $X2=1.465 $Y2=0.46
r93 2 30 150 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=4 $X=0.545
+ $Y=2.315 $X2=1.01 $Y2=2.46
r94 1 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.37 $X2=0.3 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%SCE 3 6 7 8 11 13 15 17 20 22 23 24 25 26
+ 27 34 38
c71 38 0 1.6277e-19 $X=2.395 $Y=1.295
c72 13 0 1.24551e-19 $X=1.625 $Y=2.105
r73 38 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.295
+ $X2=2.395 $Y2=1.13
r74 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=1.295 $X2=2.395 $Y2=1.295
r75 34 36 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.677 $Y=1.295
+ $X2=0.677 $Y2=1.13
r76 27 39 13.9347 $w=1.93e-07 $l=2.45e-07 $layer=LI1_cond $X=2.64 $Y=1.297
+ $X2=2.395 $Y2=1.297
r77 26 39 13.366 $w=1.93e-07 $l=2.35e-07 $layer=LI1_cond $X=2.16 $Y=1.297
+ $X2=2.395 $Y2=1.297
r78 25 26 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.297
+ $X2=2.16 $Y2=1.297
r79 24 25 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.297
+ $X2=1.68 $Y2=1.297
r80 23 24 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.297
+ $X2=1.2 $Y2=1.297
r81 23 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.295 $X2=0.75 $Y2=1.295
r82 20 40 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.485 $Y=0.615
+ $X2=2.485 $Y2=1.13
r83 15 17 110.86 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.7 $Y=2.18 $X2=1.7
+ $Y2=2.525
r84 14 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.3 $Y=2.105
+ $X2=1.225 $Y2=2.105
r85 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.625 $Y=2.105
+ $X2=1.7 $Y2=2.18
r86 13 14 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.625 $Y=2.105
+ $X2=1.3 $Y2=2.105
r87 9 22 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.225 $Y=2.18
+ $X2=1.225 $Y2=2.105
r88 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.225 $Y=2.18
+ $X2=1.225 $Y2=2.635
r89 7 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.15 $Y=2.105
+ $X2=1.225 $Y2=2.105
r90 7 8 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=1.15 $Y=2.105 $X2=0.915
+ $Y2=2.105
r91 6 8 37.7275 $w=1.5e-07 $l=2.72936e-07 $layer=POLY_cond $X=0.677 $Y=2.03
+ $X2=0.915 $Y2=2.105
r92 5 34 8.43012 $w=4.75e-07 $l=7.2e-08 $layer=POLY_cond $X=0.677 $Y=1.367
+ $X2=0.677 $Y2=1.295
r93 5 6 77.6274 $w=4.75e-07 $l=6.63e-07 $layer=POLY_cond $X=0.677 $Y=1.367
+ $X2=0.677 $Y2=2.03
r94 3 36 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.515 $Y=0.58
+ $X2=0.515 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%D 3 7 9 10 11 12 18
c35 12 0 1.24551e-19 $X=2.16 $Y=1.665
c36 7 0 8.50188e-20 $X=2.06 $Y=2.525
r37 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.655 $X2=1.825 $Y2=1.655
r38 12 19 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=2.16 $Y=1.685
+ $X2=1.825 $Y2=1.685
r39 11 19 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.685
+ $X2=1.825 $Y2=1.685
r40 10 11 23.0489 $w=2.38e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.685
+ $X2=1.68 $Y2=1.685
r41 9 10 23.0489 $w=2.38e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.685 $X2=1.2
+ $Y2=1.685
r42 5 18 38.3966 $w=2.95e-07 $l=3.1229e-07 $layer=POLY_cond $X=2.06 $Y=1.82
+ $X2=1.825 $Y2=1.64
r43 5 7 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.06 $Y=1.82 $X2=2.06
+ $Y2=2.525
r44 1 18 18.5736 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.825 $Y=1.46
+ $X2=1.825 $Y2=1.64
r45 1 3 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=1.825 $Y=1.46 $X2=1.825
+ $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%SCD 3 7 11 13 14 15 16 21
c46 3 0 3.56444e-20 $X=2.845 $Y=0.615
r47 15 16 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.137 $Y=1.665
+ $X2=3.137 $Y2=2.035
r48 14 15 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.137 $Y=1.295
+ $X2=3.137 $Y2=1.665
r49 14 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.05
+ $Y=1.34 $X2=3.05 $Y2=1.34
r50 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.05 $Y=1.68
+ $X2=3.05 $Y2=1.34
r51 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.68
+ $X2=3.05 $Y2=1.845
r52 11 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.05 $Y=1.325
+ $X2=3.05 $Y2=1.34
r53 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.992 $Y=1.175
+ $X2=2.992 $Y2=1.325
r54 7 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.96 $Y=2.525
+ $X2=2.96 $Y2=1.845
r55 3 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.845 $Y=0.615
+ $X2=2.845 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_757_317# 1 2 9 13 14 16 19 22 23 27 28
+ 32 35 36 37 38 39 40 43 52 53 56 61 62 63
c205 62 0 8.3902e-20 $X=4.9 $Y=1.29
c206 40 0 1.85618e-19 $X=7.585 $Y=1.295
c207 28 0 3.68148e-20 $X=7.955 $Y=2.22
c208 27 0 2.82467e-20 $X=7.955 $Y=2.22
c209 23 0 1.53911e-19 $X=7.77 $Y=1.26
c210 9 0 1.66968e-19 $X=3.97 $Y=2.525
r211 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.44
+ $Y=1.26 $X2=7.44 $Y2=1.26
r212 61 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=1.29
+ $X2=4.9 $Y2=1.125
r213 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.29 $X2=4.9 $Y2=1.29
r214 56 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.75
+ $X2=3.95 $Y2=1.915
r215 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.75 $X2=3.95 $Y2=1.75
r216 53 84 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=10.38 $Y=1.295
+ $X2=10.38 $Y2=2.035
r217 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=1.295
+ $X2=10.32 $Y2=1.295
r218 49 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.295
+ $X2=7.44 $Y2=1.295
r219 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r220 43 57 14.5656 $w=3.58e-07 $l=4.55e-07 $layer=LI1_cond $X=4.035 $Y=1.295
+ $X2=4.035 $Y2=1.75
r221 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.295
r222 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.295
+ $X2=7.44 $Y2=1.295
r223 39 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=10.32 $Y2=1.295
r224 39 40 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=7.585 $Y2=1.295
r225 38 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.295
+ $X2=5.04 $Y2=1.295
r226 37 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=1.295
+ $X2=7.44 $Y2=1.295
r227 37 38 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.295 $Y=1.295
+ $X2=5.185 $Y2=1.295
r228 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.295
+ $X2=4.08 $Y2=1.295
r229 35 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=5.04 $Y2=1.295
r230 35 36 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=4.225 $Y2=1.295
r231 34 53 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.38 $Y=1.165
+ $X2=10.38 $Y2=1.295
r232 32 34 2.82206 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=10.395 $Y=1.08
+ $X2=10.395 $Y2=1.165
r233 28 69 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=7.955 $Y=2.22
+ $X2=7.815 $Y2=2.22
r234 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.955
+ $Y=2.22 $X2=7.955 $Y2=2.22
r235 24 27 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=7.855 $Y=2.18
+ $X2=7.955 $Y2=2.18
r236 23 68 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=7.77 $Y=1.26
+ $X2=7.44 $Y2=1.26
r237 22 24 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.855 $Y=2.055
+ $X2=7.855 $Y2=2.18
r238 21 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.855 $Y=1.425
+ $X2=7.77 $Y2=1.26
r239 21 22 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.855 $Y=1.425
+ $X2=7.855 $Y2=2.055
r240 17 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.815 $Y=2.385
+ $X2=7.815 $Y2=2.22
r241 17 19 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.815 $Y=2.385
+ $X2=7.815 $Y2=2.875
r242 14 67 53.3511 $w=2.62e-07 $l=3.63249e-07 $layer=POLY_cond $X=7.15 $Y=1.095
+ $X2=7.44 $Y2=1.26
r243 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.15 $Y=1.095
+ $X2=7.15 $Y2=0.775
r244 13 63 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.88 $Y=0.805
+ $X2=4.88 $Y2=1.125
r245 9 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.97 $Y=2.525
+ $X2=3.97 $Y2=1.915
r246 2 84 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=10.28
+ $Y=1.835 $X2=10.405 $Y2=2.035
r247 1 32 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=10.265
+ $Y=0.785 $X2=10.41 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_937_333# 1 2 9 11 15 18 20 21 25 28 29
+ 31 33 39 43
c98 39 0 2.9296e-19 $X=6.74 $Y=1.685
c99 33 0 1.16283e-19 $X=4.87 $Y=1.685
c100 31 0 5.31087e-20 $X=6.98 $Y=2.055
c101 28 0 1.85378e-20 $X=6.745 $Y=1.96
c102 21 0 7.65474e-20 $X=6.645 $Y=1.685
r103 37 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.83
+ $X2=5.015 $Y2=1.83
r104 37 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.85 $Y=1.83 $X2=4.76
+ $Y2=1.83
r105 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.83 $X2=4.85 $Y2=1.83
r106 33 36 5.76222 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=4.87 $Y=1.685
+ $X2=4.87 $Y2=1.83
r107 29 31 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=6.835 $Y=2.055
+ $X2=6.98 $Y2=2.055
r108 28 29 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=6.745 $Y=1.96
+ $X2=6.835 $Y2=2.055
r109 27 39 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.745 $Y=1.77
+ $X2=6.74 $Y2=1.685
r110 27 28 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=6.745 $Y=1.77
+ $X2=6.745 $Y2=1.96
r111 23 39 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.74 $Y=1.6
+ $X2=6.74 $Y2=1.685
r112 23 25 46.9904 $w=1.88e-07 $l=8.05e-07 $layer=LI1_cond $X=6.74 $Y=1.6
+ $X2=6.74 $Y2=0.795
r113 22 33 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.015 $Y=1.685
+ $X2=4.87 $Y2=1.685
r114 21 39 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.645 $Y=1.685
+ $X2=6.74 $Y2=1.685
r115 21 22 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=6.645 $Y=1.685
+ $X2=5.015 $Y2=1.685
r116 19 20 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.365 $Y=1.275
+ $X2=5.365 $Y2=1.425
r117 18 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.38 $Y=1.695
+ $X2=5.38 $Y2=1.425
r118 15 19 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.35 $Y=0.805 $X2=5.35
+ $Y2=1.275
r119 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.305 $Y=1.77
+ $X2=5.38 $Y2=1.695
r120 11 43 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.305 $Y=1.77
+ $X2=5.015 $Y2=1.77
r121 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.76 $Y=1.995
+ $X2=4.76 $Y2=1.83
r122 7 9 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.76 $Y=1.995
+ $X2=4.76 $Y2=2.525
r123 2 31 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.895 $X2=6.98 $Y2=2.055
r124 1 25 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=6.6
+ $Y=0.565 $X2=6.74 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%RESET_B 3 5 6 11 12 13 15 16 18 20 21 22
+ 28 31 35 37 38 39 41 42 45 46 47 49 50 51 53 56 57 62 64 70
c207 70 0 6.31513e-20 $X=9.24 $Y=2.34
c208 41 0 1.60449e-19 $X=5.845 $Y=1.245
c209 31 0 2.92081e-20 $X=9.015 $Y=0.805
c210 16 0 1.14005e-19 $X=5.785 $Y=0.18
c211 15 0 5.71712e-20 $X=3.845 $Y=1.195
c212 12 0 9.02003e-20 $X=3.77 $Y=1.27
r213 62 64 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=5.942 $Y=2.04
+ $X2=5.942 $Y2=1.875
r214 56 57 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=5.965 $Y=2.035
+ $X2=5.965 $Y2=2.32
r215 56 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.965
+ $Y=2.04 $X2=5.965 $Y2=2.04
r216 54 70 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=9.105 $Y=2.34
+ $X2=9.24 $Y2=2.34
r217 54 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.105 $Y=2.34
+ $X2=9.015 $Y2=2.34
r218 53 55 8.41379 $w=3.19e-07 $l=2.2e-07 $layer=LI1_cond $X=9.105 $Y=2.34
+ $X2=9.105 $Y2=2.56
r219 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.105
+ $Y=2.34 $X2=9.105 $Y2=2.34
r220 50 55 4.42298 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.94 $Y=2.56
+ $X2=9.105 $Y2=2.56
r221 50 51 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.94 $Y=2.56
+ $X2=8.285 $Y2=2.56
r222 48 51 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.16 $Y=2.645
+ $X2=8.285 $Y2=2.56
r223 48 49 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=8.16 $Y=2.645
+ $X2=8.16 $Y2=2.905
r224 46 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.035 $Y=2.99
+ $X2=8.16 $Y2=2.905
r225 46 47 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=8.035 $Y=2.99
+ $X2=6.95 $Y2=2.99
r226 45 47 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.86 $Y=2.905
+ $X2=6.95 $Y2=2.99
r227 44 45 25.5707 $w=1.78e-07 $l=4.15e-07 $layer=LI1_cond $X=6.86 $Y=2.49
+ $X2=6.86 $Y2=2.905
r228 43 57 4.90495 $w=1.7e-07 $l=1.77989e-07 $layer=LI1_cond $X=6.13 $Y=2.405
+ $X2=5.965 $Y2=2.432
r229 42 44 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.77 $Y=2.405
+ $X2=6.86 $Y2=2.49
r230 42 43 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.77 $Y=2.405
+ $X2=6.13 $Y2=2.405
r231 41 64 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=5.83 $Y=1.245
+ $X2=5.83 $Y2=1.875
r232 40 41 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.845 $Y=1.095
+ $X2=5.845 $Y2=1.245
r233 37 38 41.3657 $w=1.9e-07 $l=1.15e-07 $layer=POLY_cond $X=3.52 $Y=2.125
+ $X2=3.52 $Y2=2.24
r234 33 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.24 $Y=2.505
+ $X2=9.24 $Y2=2.34
r235 33 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.24 $Y=2.505
+ $X2=9.24 $Y2=2.875
r236 29 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.015 $Y=2.175
+ $X2=9.015 $Y2=2.34
r237 29 31 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=9.015 $Y=2.175
+ $X2=9.015 $Y2=0.805
r238 28 40 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.86 $Y=0.775
+ $X2=5.86 $Y2=1.095
r239 25 28 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.86 $Y=0.255
+ $X2=5.86 $Y2=0.775
r240 21 62 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=5.942 $Y=2.13
+ $X2=5.942 $Y2=2.04
r241 21 22 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=5.755 $Y=2.13
+ $X2=5.375 $Y2=2.13
r242 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.3 $Y=2.205
+ $X2=5.375 $Y2=2.13
r243 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.3 $Y=2.205
+ $X2=5.3 $Y2=2.525
r244 17 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.92 $Y=0.18
+ $X2=3.845 $Y2=0.18
r245 16 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=5.86 $Y2=0.255
r246 16 17 956.309 $w=1.5e-07 $l=1.865e-06 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=3.92 $Y2=0.18
r247 14 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.845 $Y=0.255
+ $X2=3.845 $Y2=0.18
r248 14 15 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.845 $Y=0.255
+ $X2=3.845 $Y2=1.195
r249 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.77 $Y=1.27
+ $X2=3.845 $Y2=1.195
r250 12 13 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.77 $Y=1.27
+ $X2=3.575 $Y2=1.27
r251 11 38 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.54 $Y=2.525
+ $X2=3.54 $Y2=2.24
r252 7 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=1.345
+ $X2=3.575 $Y2=1.27
r253 7 37 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.5 $Y=1.345 $X2=3.5
+ $Y2=2.125
r254 5 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=0.18
+ $X2=3.845 $Y2=0.18
r255 5 6 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=3.77 $Y=0.18
+ $X2=3.395 $Y2=0.18
r256 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.32 $Y=0.255
+ $X2=3.395 $Y2=0.18
r257 1 3 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.32 $Y=0.255
+ $X2=3.32 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_809_463# 1 2 3 12 14 16 19 22 23 24 27
+ 31 34 35 37 43 45
c124 43 0 8.63327e-20 $X=4.555 $Y=2.21
c125 24 0 5.71712e-20 $X=4.555 $Y=0.89
c126 23 0 1.16283e-19 $X=5.465 $Y=0.89
c127 14 0 5.31087e-20 $X=6.765 $Y=1.635
r128 42 43 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.47 $Y=2.21
+ $X2=4.555 $Y2=2.21
r129 38 45 29.1096 $w=3.56e-07 $l=2.15e-07 $layer=POLY_cond $X=6.31 $Y=1.402
+ $X2=6.525 $Y2=1.402
r130 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=1.335 $X2=6.31 $Y2=1.335
r131 35 37 28.3678 $w=2.58e-07 $l=6.4e-07 $layer=LI1_cond $X=5.67 $Y=1.3
+ $X2=6.31 $Y2=1.3
r132 34 35 6.94126 $w=2.6e-07 $l=1.7404e-07 $layer=LI1_cond $X=5.567 $Y=1.17
+ $X2=5.67 $Y2=1.3
r133 33 34 9.46785 $w=2.03e-07 $l=1.75e-07 $layer=LI1_cond $X=5.567 $Y=0.995
+ $X2=5.567 $Y2=1.17
r134 29 31 8.2628 $w=2.63e-07 $l=1.9e-07 $layer=LI1_cond $X=5.497 $Y=2.335
+ $X2=5.497 $Y2=2.525
r135 27 29 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.365 $Y=2.25
+ $X2=5.497 $Y2=2.335
r136 27 43 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.365 $Y=2.25
+ $X2=4.555 $Y2=2.25
r137 24 26 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=4.555 $Y=0.89
+ $X2=4.665 $Y2=0.89
r138 23 33 6.81778 $w=2.1e-07 $l=1.47428e-07 $layer=LI1_cond $X=5.465 $Y=0.89
+ $X2=5.567 $Y2=0.995
r139 23 26 42.2511 $w=2.08e-07 $l=8e-07 $layer=LI1_cond $X=5.465 $Y=0.89
+ $X2=4.665 $Y2=0.89
r140 22 42 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.47 $Y=2.085
+ $X2=4.47 $Y2=2.21
r141 21 24 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.47 $Y=0.995
+ $X2=4.555 $Y2=0.89
r142 21 22 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=2.085
r143 17 42 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=4.225 $Y=2.21
+ $X2=4.47 $Y2=2.21
r144 17 19 6.84263 $w=3.18e-07 $l=1.9e-07 $layer=LI1_cond $X=4.225 $Y=2.335
+ $X2=4.225 $Y2=2.525
r145 14 45 32.4944 $w=3.56e-07 $l=3.36927e-07 $layer=POLY_cond $X=6.765 $Y=1.635
+ $X2=6.525 $Y2=1.402
r146 14 16 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=6.765 $Y=1.635
+ $X2=6.765 $Y2=2.105
r147 10 45 23.0368 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=1.402
r148 10 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=0.775
r149 3 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=2.315 $X2=5.515 $Y2=2.525
r150 2 19 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=2.315 $X2=4.185 $Y2=2.525
r151 1 26 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.595 $X2=4.665 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_865_255# 1 2 10 13 15 16 20 21 22 25 27
+ 29 30 32 34 36 37 40 41 42 44 48 51 53 55 57 58 62 67 72
c208 72 0 6.71069e-20 $X=10.625 $Y=1.51
c209 55 0 1.23014e-19 $X=10.8 $Y=1.51
c210 53 0 2.24062e-19 $X=8.37 $Y=1.65
c211 36 0 1.80416e-19 $X=7.815 $Y=1.635
c212 34 0 8.63327e-20 $X=4.425 $Y=1.425
c213 22 0 1.54882e-19 $X=7.27 $Y=1.71
c214 21 0 2.82467e-20 $X=7.815 $Y=1.71
r215 71 72 0.734756 $w=3.28e-07 $l=5e-09 $layer=POLY_cond $X=10.62 $Y=1.51
+ $X2=10.625 $Y2=1.51
r216 64 67 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=11.295 $Y=2.88
+ $X2=11.465 $Y2=2.88
r217 59 62 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=11.29 $Y=1.085
+ $X2=11.465 $Y2=1.085
r218 56 72 25.7165 $w=3.28e-07 $l=1.75e-07 $layer=POLY_cond $X=10.8 $Y=1.51
+ $X2=10.625 $Y2=1.51
r219 55 57 10.1645 $w=6.63e-07 $l=1.65e-07 $layer=LI1_cond $X=11.047 $Y=1.51
+ $X2=11.047 $Y2=1.345
r220 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.8
+ $Y=1.51 $X2=10.8 $Y2=1.51
r221 50 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=1.65
+ $X2=8.37 $Y2=1.65
r222 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.205
+ $Y=1.65 $X2=8.205 $Y2=1.65
r223 48 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.295 $Y=2.715
+ $X2=11.295 $Y2=2.88
r224 47 58 2.32396 $w=4.17e-07 $l=2.87374e-07 $layer=LI1_cond $X=11.295 $Y=2.54
+ $X2=11.047 $Y2=2.455
r225 47 48 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=11.295 $Y=2.54
+ $X2=11.295 $Y2=2.715
r226 45 59 1.35108 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=11.29 $Y=1.185
+ $X2=11.29 $Y2=1.085
r227 45 57 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=11.29 $Y=1.185
+ $X2=11.29 $Y2=1.345
r228 44 58 2.32396 $w=4.17e-07 $l=8.5e-08 $layer=LI1_cond $X=11.047 $Y=2.37
+ $X2=11.047 $Y2=2.455
r229 43 55 3.00369 $w=6.63e-07 $l=1.67e-07 $layer=LI1_cond $X=11.047 $Y=1.677
+ $X2=11.047 $Y2=1.51
r230 43 44 12.4644 $w=6.63e-07 $l=6.93e-07 $layer=LI1_cond $X=11.047 $Y=1.677
+ $X2=11.047 $Y2=2.37
r231 41 58 4.70729 $w=1.7e-07 $l=3.32e-07 $layer=LI1_cond $X=10.715 $Y=2.455
+ $X2=11.047 $Y2=2.455
r232 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.715 $Y=2.455
+ $X2=10.045 $Y2=2.455
r233 40 42 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=9.922 $Y=2.37
+ $X2=10.045 $Y2=2.455
r234 39 40 30.3398 $w=2.43e-07 $l=6.45e-07 $layer=LI1_cond $X=9.922 $Y=1.725
+ $X2=9.922 $Y2=2.37
r235 37 39 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=9.8 $Y=1.64
+ $X2=9.922 $Y2=1.725
r236 37 53 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=9.8 $Y=1.64
+ $X2=8.37 $Y2=1.64
r237 35 51 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.995 $Y=1.65
+ $X2=8.205 $Y2=1.65
r238 35 36 13.5877 $w=2.4e-07 $l=1.8735e-07 $layer=POLY_cond $X=7.995 $Y=1.65
+ $X2=7.815 $Y2=1.635
r239 33 34 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.425 $Y=1.275
+ $X2=4.425 $Y2=1.425
r240 30 72 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.625 $Y=1.345
+ $X2=10.625 $Y2=1.51
r241 30 32 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=10.625 $Y=1.345
+ $X2=10.625 $Y2=0.995
r242 27 71 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.62 $Y=1.675
+ $X2=10.62 $Y2=1.51
r243 27 29 118.893 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.62 $Y=1.675
+ $X2=10.62 $Y2=2.045
r244 23 36 12.1617 $w=1.5e-07 $l=1.95576e-07 $layer=POLY_cond $X=7.92 $Y=1.485
+ $X2=7.815 $Y2=1.635
r245 23 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.92 $Y=1.485
+ $X2=7.92 $Y2=0.775
r246 21 36 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=7.815 $Y=1.71
+ $X2=7.815 $Y2=1.635
r247 21 22 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.815 $Y=1.71
+ $X2=7.27 $Y2=1.71
r248 18 20 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.195 $Y=3.075
+ $X2=7.195 $Y2=2.105
r249 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.195 $Y=1.785
+ $X2=7.27 $Y2=1.71
r250 17 20 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.195 $Y=1.785
+ $X2=7.195 $Y2=2.105
r251 15 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.12 $Y=3.15
+ $X2=7.195 $Y2=3.075
r252 15 16 1356.27 $w=1.5e-07 $l=2.645e-06 $layer=POLY_cond $X=7.12 $Y=3.15
+ $X2=4.475 $Y2=3.15
r253 13 33 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.45 $Y=0.805 $X2=4.45
+ $Y2=1.275
r254 10 34 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=4.4 $Y=2.525
+ $X2=4.4 $Y2=1.425
r255 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.4 $Y=3.075
+ $X2=4.475 $Y2=3.15
r256 8 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.4 $Y=3.075 $X2=4.4
+ $Y2=2.525
r257 2 67 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=11.325
+ $Y=2.675 $X2=11.465 $Y2=2.88
r258 1 62 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=11.325
+ $Y=0.785 $X2=11.465 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_1445_113# 1 2 7 9 12 16 20 24 26 28 29
+ 31 35 36 39 42 44 46 47 48 50 58 61 62 63 68 69
c207 68 0 3.17486e-19 $X=12.29 $Y=1.08
c208 44 0 1.85618e-19 $X=8.32 $Y=1.22
c209 31 0 9.19974e-20 $X=7.41 $Y=2.04
c210 29 0 8.84191e-20 $X=7.445 $Y=1.79
r211 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.29
+ $Y=1.08 $X2=12.29 $Y2=1.08
r212 65 68 24.3384 $w=1.78e-07 $l=3.95e-07 $layer=LI1_cond $X=11.895 $Y=1.075
+ $X2=12.29 $Y2=1.075
r213 61 74 4.53008 $w=2.66e-07 $l=2.5e-08 $layer=POLY_cond $X=9.645 $Y=1.29
+ $X2=9.67 $Y2=1.29
r214 60 63 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=9.645 $Y=1.26
+ $X2=9.96 $Y2=1.26
r215 60 62 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.645 $Y=1.26
+ $X2=9.48 $Y2=1.26
r216 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.645
+ $Y=1.29 $X2=9.645 $Y2=1.29
r217 50 65 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=11.895 $Y=0.985
+ $X2=11.895 $Y2=1.075
r218 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.895 $Y=0.815
+ $X2=11.895 $Y2=0.985
r219 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.81 $Y=0.73
+ $X2=11.895 $Y2=0.815
r220 47 48 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=11.81 $Y=0.73
+ $X2=10.045 $Y2=0.73
r221 46 63 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.96 $Y=1.135
+ $X2=9.96 $Y2=1.26
r222 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.96 $Y=0.815
+ $X2=10.045 $Y2=0.73
r223 45 46 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.96 $Y=0.815
+ $X2=9.96 $Y2=1.135
r224 44 62 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=8.32 $Y=1.22
+ $X2=9.48 $Y2=1.22
r225 42 44 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.215 $Y=1.135
+ $X2=8.32 $Y2=1.22
r226 41 42 11.619 $w=2.08e-07 $l=2.2e-07 $layer=LI1_cond $X=8.215 $Y=0.915
+ $X2=8.215 $Y2=1.135
r227 39 41 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.11 $Y=0.83
+ $X2=8.215 $Y2=0.915
r228 39 58 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.11 $Y=0.83
+ $X2=7.87 $Y2=0.83
r229 36 53 11.4481 $w=2.9e-07 $l=2.55e-07 $layer=LI1_cond $X=7.345 $Y=0.77
+ $X2=7.09 $Y2=0.77
r230 36 38 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.345 $Y=0.77
+ $X2=7.705 $Y2=0.77
r231 35 58 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=7.725 $Y=0.77
+ $X2=7.87 $Y2=0.77
r232 35 38 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=7.725 $Y=0.77
+ $X2=7.705 $Y2=0.77
r233 31 33 23.4921 $w=2.58e-07 $l=5.3e-07 $layer=LI1_cond $X=7.445 $Y=2.04
+ $X2=7.445 $Y2=2.57
r234 29 54 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.445 $Y=1.705
+ $X2=7.09 $Y2=1.705
r235 29 31 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=7.445 $Y=1.79
+ $X2=7.445 $Y2=2.04
r236 28 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.62
+ $X2=7.09 $Y2=1.705
r237 27 53 2.27611 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.09 $Y=0.915
+ $X2=7.09 $Y2=0.77
r238 27 28 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.09 $Y=0.915
+ $X2=7.09 $Y2=1.62
r239 25 69 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=12.29 $Y=1.42
+ $X2=12.29 $Y2=1.08
r240 25 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.29 $Y=1.42
+ $X2=12.29 $Y2=1.585
r241 24 69 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=12.29 $Y=1.065
+ $X2=12.29 $Y2=1.08
r242 23 24 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=12.327 $Y=0.915
+ $X2=12.327 $Y2=1.065
r243 20 23 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=12.455 $Y=0.445
+ $X2=12.455 $Y2=0.915
r244 16 26 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=12.38 $Y=2.155
+ $X2=12.38 $Y2=1.585
r245 10 74 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.67 $Y=1.455
+ $X2=9.67 $Y2=1.29
r246 10 12 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=9.67 $Y=1.455
+ $X2=9.67 $Y2=2.875
r247 7 61 48.9248 $w=2.66e-07 $l=3.4271e-07 $layer=POLY_cond $X=9.375 $Y=1.125
+ $X2=9.645 $Y2=1.29
r248 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.375 $Y=1.125
+ $X2=9.375 $Y2=0.805
r249 2 33 600 $w=1.7e-07 $l=7.68521e-07 $layer=licon1_PDIFF $count=1 $X=7.27
+ $Y=1.895 $X2=7.47 $Y2=2.57
r250 2 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.27
+ $Y=1.895 $X2=7.41 $Y2=2.04
r251 1 38 91 $w=1.7e-07 $l=5.81722e-07 $layer=licon1_NDIFF $count=2 $X=7.225
+ $Y=0.565 $X2=7.705 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_1641_21# 1 2 10 13 15 16 17 18 20 21 25
+ 29 31 34 39 40 45 47
c113 34 0 6.31513e-20 $X=8.565 $Y=1.99
c114 29 0 2.92081e-20 $X=9.705 $Y=0.365
c115 18 0 3.41158e-19 $X=8.355 $Y=1.17
r116 39 40 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.49 $Y=2.91
+ $X2=9.49 $Y2=2.745
r117 37 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.565 $Y=2.22
+ $X2=8.655 $Y2=2.22
r118 37 42 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=8.565 $Y=2.22
+ $X2=8.405 $Y2=2.22
r119 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.565
+ $Y=2.22 $X2=8.565 $Y2=2.22
r120 34 36 10.3926 $w=2.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.565 $Y=1.99
+ $X2=8.565 $Y2=2.22
r121 32 47 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=9.99 $Y=0.35
+ $X2=9.99 $Y2=0.18
r122 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.99
+ $Y=0.35 $X2=9.99 $Y2=0.35
r123 29 31 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=9.705 $Y=0.365
+ $X2=9.99 $Y2=0.365
r124 27 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.535 $Y=2.075
+ $X2=9.535 $Y2=2.745
r125 23 29 6.94494 $w=2.2e-07 $l=1.87083e-07 $layer=LI1_cond $X=9.565 $Y=0.475
+ $X2=9.705 $Y2=0.365
r126 23 25 13.3766 $w=2.78e-07 $l=3.25e-07 $layer=LI1_cond $X=9.565 $Y=0.475
+ $X2=9.565 $Y2=0.8
r127 22 34 3.44395 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.73 $Y=1.99
+ $X2=8.565 $Y2=1.99
r128 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.45 $Y=1.99
+ $X2=9.535 $Y2=2.075
r129 21 22 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=9.45 $Y=1.99
+ $X2=8.73 $Y2=1.99
r130 20 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=2.055
+ $X2=8.655 $Y2=2.22
r131 19 20 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=8.655 $Y=1.245
+ $X2=8.655 $Y2=2.055
r132 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.58 $Y=1.17
+ $X2=8.655 $Y2=1.245
r133 17 18 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=8.58 $Y=1.17
+ $X2=8.355 $Y2=1.17
r134 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.825 $Y=0.18
+ $X2=9.99 $Y2=0.18
r135 15 16 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=9.825 $Y=0.18
+ $X2=8.355 $Y2=0.18
r136 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.405 $Y=2.385
+ $X2=8.405 $Y2=2.22
r137 11 13 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.405 $Y=2.385
+ $X2=8.405 $Y2=2.875
r138 8 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.28 $Y=1.095
+ $X2=8.355 $Y2=1.17
r139 8 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.28 $Y=1.095
+ $X2=8.28 $Y2=0.775
r140 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.28 $Y=0.255
+ $X2=8.355 $Y2=0.18
r141 7 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.28 $Y=0.255
+ $X2=8.28 $Y2=0.775
r142 2 39 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=9.315
+ $Y=2.665 $X2=9.455 $Y2=2.91
r143 1 25 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=9.45
+ $Y=0.595 $X2=9.59 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%CLK 1 3 6 8 10 11 12 13 17 21
c46 21 0 2.35015e-19 $X=11.715 $Y=1.51
r47 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.715
+ $Y=1.51 $X2=11.715 $Y2=1.51
r48 17 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.715 $Y=1.42
+ $X2=11.715 $Y2=1.51
r49 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.715 $Y=2.035
+ $X2=11.715 $Y2=2.405
r50 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.715 $Y=1.665
+ $X2=11.715 $Y2=2.035
r51 11 21 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=11.715 $Y=1.665
+ $X2=11.715 $Y2=1.51
r52 9 10 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.325 $Y=1.42
+ $X2=11.25 $Y2=1.42
r53 8 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.55 $Y=1.42
+ $X2=11.715 $Y2=1.42
r54 8 9 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=11.55 $Y=1.42
+ $X2=11.325 $Y2=1.42
r55 4 10 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.25 $Y=1.495
+ $X2=11.25 $Y2=1.42
r56 4 6 712.745 $w=1.5e-07 $l=1.39e-06 $layer=POLY_cond $X=11.25 $Y=1.495
+ $X2=11.25 $Y2=2.885
r57 1 10 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.25 $Y=1.345
+ $X2=11.25 $Y2=1.42
r58 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11.25 $Y=1.345
+ $X2=11.25 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_2408_367# 1 2 9 13 17 21 23 24 25 26 30
+ 31
c57 30 0 1.96847e-19 $X=12.83 $Y=1.47
c58 23 0 2.77631e-20 $X=12.665 $Y=1.76
c59 9 0 2.89723e-19 $X=12.965 $Y=0.655
r60 31 34 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.852 $Y=1.47
+ $X2=12.852 $Y2=1.635
r61 31 33 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.852 $Y=1.47
+ $X2=12.852 $Y2=1.305
r62 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.83
+ $Y=1.47 $X2=12.83 $Y2=1.47
r63 28 30 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=12.79 $Y=1.675
+ $X2=12.79 $Y2=1.47
r64 27 30 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=12.79 $Y=0.815
+ $X2=12.79 $Y2=1.47
r65 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.665 $Y=0.73
+ $X2=12.79 $Y2=0.815
r66 25 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.665 $Y=0.73
+ $X2=12.405 $Y2=0.73
r67 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.665 $Y=1.76
+ $X2=12.79 $Y2=1.675
r68 23 24 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=12.665 $Y=1.76
+ $X2=12.26 $Y2=1.76
r69 19 26 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=12.277 $Y=0.645
+ $X2=12.405 $Y2=0.73
r70 19 21 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=12.277 $Y=0.645
+ $X2=12.277 $Y2=0.44
r71 15 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=12.155 $Y=1.845
+ $X2=12.26 $Y2=1.76
r72 15 17 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=12.155 $Y=1.845
+ $X2=12.155 $Y2=1.98
r73 13 34 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=12.965 $Y=2.465
+ $X2=12.965 $Y2=1.635
r74 9 33 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=12.965 $Y=0.655
+ $X2=12.965 $Y2=1.305
r75 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.04
+ $Y=1.835 $X2=12.165 $Y2=1.98
r76 1 21 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=12.115
+ $Y=0.235 $X2=12.24 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 41 45 47
+ 51 55 60 61 62 71 75 83 96 106 107 110 113 116 121 124 126 129 132
c150 55 0 1.67908e-19 $X=12.595 $Y=2.1
r151 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r152 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r153 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r154 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r155 123 124 9.89636 $w=5.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=3.135
+ $X2=9.19 $Y2=3.135
r156 120 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r157 119 123 3.09699 $w=5.58e-07 $l=1.45e-07 $layer=LI1_cond $X=8.88 $Y=3.135
+ $X2=9.025 $Y2=3.135
r158 119 121 15.4496 $w=5.58e-07 $l=4.25e-07 $layer=LI1_cond $X=8.88 $Y=3.135
+ $X2=8.455 $Y2=3.135
r159 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r160 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r161 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r162 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r163 107 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r164 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r165 104 132 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=12.915 $Y=3.33
+ $X2=12.672 $Y2=3.33
r166 104 106 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.915 $Y=3.33
+ $X2=13.2 $Y2=3.33
r167 103 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r168 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r169 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r170 100 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r171 99 102 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r172 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r173 97 129 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=10.897 $Y2=3.33
r174 97 99 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=11.28 $Y2=3.33
r175 96 132 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=12.43 $Y=3.33
+ $X2=12.672 $Y2=3.33
r176 96 102 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.43 $Y=3.33
+ $X2=12.24 $Y2=3.33
r177 95 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r178 94 121 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=8.455 $Y2=3.33
r179 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r180 92 95 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r181 91 94 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r182 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r183 89 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.435 $Y2=3.33
r184 89 91 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r185 87 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r186 87 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r187 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r188 84 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=3.33
+ $X2=5.03 $Y2=3.33
r189 84 86 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=5.195 $Y=3.33
+ $X2=6 $Y2=3.33
r190 83 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.27 $Y=3.33
+ $X2=6.435 $Y2=3.33
r191 83 86 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.27 $Y=3.33 $X2=6
+ $Y2=3.33
r192 82 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r193 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r194 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r195 79 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r196 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r197 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r198 76 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=3.33
+ $X2=3.235 $Y2=3.33
r199 76 78 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r200 75 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=5.03 $Y2=3.33
r201 75 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=4.56 $Y2=3.33
r202 74 111 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r203 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r204 71 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=3.235 $Y2=3.33
r205 71 73 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=1.68 $Y2=3.33
r206 70 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r207 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r208 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r209 65 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r210 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r211 62 92 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r212 62 117 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r213 60 69 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.2 $Y2=3.33
r214 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.485 $Y2=3.33
r215 59 73 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.65 $Y=3.33 $X2=1.68
+ $Y2=3.33
r216 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.485 $Y2=3.33
r217 55 58 9.98787 $w=4.83e-07 $l=4.05e-07 $layer=LI1_cond $X=12.672 $Y=2.1
+ $X2=12.672 $Y2=2.505
r218 53 132 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=12.672 $Y=3.245
+ $X2=12.672 $Y2=3.33
r219 53 58 18.2494 $w=4.83e-07 $l=7.4e-07 $layer=LI1_cond $X=12.672 $Y=3.245
+ $X2=12.672 $Y2=2.505
r220 49 129 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=10.897 $Y=3.245
+ $X2=10.897 $Y2=3.33
r221 49 51 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=10.897 $Y=3.245
+ $X2=10.897 $Y2=2.875
r222 48 126 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.05 $Y=3.33
+ $X2=9.92 $Y2=3.33
r223 47 129 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=10.755 $Y=3.33
+ $X2=10.897 $Y2=3.33
r224 47 48 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=10.755 $Y=3.33
+ $X2=10.05 $Y2=3.33
r225 43 126 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.92 $Y=3.245
+ $X2=9.92 $Y2=3.33
r226 43 45 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=9.92 $Y=3.245
+ $X2=9.92 $Y2=2.875
r227 41 126 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.79 $Y=3.33
+ $X2=9.92 $Y2=3.33
r228 41 124 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=9.79 $Y=3.33
+ $X2=9.19 $Y2=3.33
r229 37 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=3.245
+ $X2=6.435 $Y2=3.33
r230 37 39 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.435 $Y=3.245
+ $X2=6.435 $Y2=2.755
r231 33 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=3.33
r232 33 35 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=2.61
r233 29 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=3.245
+ $X2=3.235 $Y2=3.33
r234 29 31 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.235 $Y=3.245
+ $X2=3.235 $Y2=2.77
r235 25 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=3.33
r236 25 27 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=2.555
r237 8 58 300 $w=1.7e-07 $l=8.04083e-07 $layer=licon1_PDIFF $count=2 $X=12.455
+ $Y=1.835 $X2=12.75 $Y2=2.505
r238 8 55 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=12.455
+ $Y=1.835 $X2=12.595 $Y2=2.1
r239 7 51 600 $w=1.7e-07 $l=1.147e-06 $layer=licon1_PDIFF $count=1 $X=10.695
+ $Y=1.835 $X2=10.92 $Y2=2.875
r240 6 45 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.745
+ $Y=2.665 $X2=9.885 $Y2=2.875
r241 5 123 300 $w=1.7e-07 $l=6.76609e-07 $layer=licon1_PDIFF $count=2 $X=8.48
+ $Y=2.665 $X2=9.025 $Y2=2.96
r242 4 39 600 $w=1.7e-07 $l=9.29677e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.895 $X2=6.435 $Y2=2.755
r243 3 35 600 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_PDIFF $count=1 $X=4.835
+ $Y=2.315 $X2=5.03 $Y2=2.61
r244 2 31 600 $w=1.7e-07 $l=5.45917e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=2.315 $X2=3.235 $Y2=2.77
r245 1 27 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=1.3
+ $Y=2.315 $X2=1.485 $Y2=2.555
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%A_380_50# 1 2 3 4 13 15 18 19 22 26 31 32
+ 36
c94 32 0 1.66968e-19 $X=3.582 $Y=2.46
c95 31 0 8.87678e-20 $X=3.582 $Y=0.9
c96 19 0 2.10427e-19 $X=4.015 $Y=0.9
c97 15 0 2.81154e-21 $X=3.48 $Y=2.4
r98 36 38 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=4.115 $Y=0.82
+ $X2=4.115 $Y2=0.9
r99 32 34 7.25292 $w=2.91e-07 $l=1.73e-07 $layer=LI1_cond $X=3.582 $Y=2.46
+ $X2=3.755 $Y2=2.46
r100 26 29 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.275 $Y=2.4
+ $X2=2.275 $Y2=2.515
r101 22 24 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.155 $Y=0.7 $X2=2.155
+ $Y2=0.9
r102 20 31 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=3.685 $Y=0.9
+ $X2=3.582 $Y2=0.9
r103 19 38 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.015 $Y=0.9 $X2=4.115
+ $Y2=0.9
r104 19 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.015 $Y=0.9
+ $X2=3.685 $Y2=0.9
r105 18 32 2.81016 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=3.582 $Y=2.295
+ $X2=3.582 $Y2=2.46
r106 17 31 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.582 $Y=0.985
+ $X2=3.582 $Y2=0.9
r107 17 18 70.8736 $w=2.03e-07 $l=1.31e-06 $layer=LI1_cond $X=3.582 $Y=0.985
+ $X2=3.582 $Y2=2.295
r108 16 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=2.4
+ $X2=2.275 $Y2=2.4
r109 15 32 6.36801 $w=2.91e-07 $l=1.28546e-07 $layer=LI1_cond $X=3.48 $Y=2.4
+ $X2=3.582 $Y2=2.46
r110 15 16 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.48 $Y=2.4
+ $X2=2.44 $Y2=2.4
r111 14 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=0.9
+ $X2=2.155 $Y2=0.9
r112 13 31 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=3.48 $Y=0.9
+ $X2=3.582 $Y2=0.9
r113 13 14 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.48 $Y=0.9
+ $X2=2.32 $Y2=0.9
r114 4 34 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=2.315 $X2=3.755 $Y2=2.46
r115 3 29 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=2.315 $X2=2.275 $Y2=2.515
r116 2 36 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.595 $X2=4.13 $Y2=0.82
r117 1 22 182 $w=1.7e-07 $l=5.6325e-07 $layer=licon1_NDIFF $count=1 $X=1.9
+ $Y=0.25 $X2=2.155 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%Q 1 2 7 8 9 10 11 12 20
r11 12 36 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=13.22 $Y=2.775
+ $X2=13.22 $Y2=2.91
r12 11 12 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.22 $Y=2.405
+ $X2=13.22 $Y2=2.775
r13 10 11 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=13.22 $Y=1.98
+ $X2=13.22 $Y2=2.405
r14 9 10 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.22 $Y=1.665
+ $X2=13.22 $Y2=1.98
r15 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.22 $Y=1.295
+ $X2=13.22 $Y2=1.665
r16 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.22 $Y=0.925
+ $X2=13.22 $Y2=1.295
r17 7 20 21.555 $w=2.68e-07 $l=5.05e-07 $layer=LI1_cond $X=13.22 $Y=0.925
+ $X2=13.22 $Y2=0.42
r18 2 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.04
+ $Y=1.835 $X2=13.18 $Y2=2.91
r19 2 10 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.04
+ $Y=1.835 $X2=13.18 $Y2=1.98
r20 1 20 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=13.04
+ $Y=0.235 $X2=13.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45
+ 47 48 49 51 56 77 81 91 92 95 98 101 104
c140 92 0 5.91316e-20 $X=13.2 $Y=0
c141 56 0 1.18827e-19 $X=3.405 $Y=0
c142 25 0 9.02003e-20 $X=3.57 $Y=0.55
c143 2 0 9.64219e-20 $X=3.395 $Y=0.405
r144 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r145 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r146 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r147 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r148 92 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r149 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r150 89 104 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=12.745 $Y2=0
r151 89 91 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=13.2 $Y2=0
r152 88 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r153 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r154 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r155 85 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r156 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=0 $X2=12.24
+ $Y2=0
r157 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r158 82 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.92 $Y2=0
r159 82 84 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.28 $Y2=0
r160 81 104 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.575 $Y=0
+ $X2=12.745 $Y2=0
r161 81 87 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.575 $Y=0
+ $X2=12.24 $Y2=0
r162 80 102 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.8 $Y2=0
r163 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r164 77 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=10.92 $Y2=0
r165 77 79 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=8.88 $Y2=0
r166 76 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r167 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r168 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r169 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r170 70 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r171 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r172 67 70 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r173 67 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r174 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r175 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r176 64 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.57
+ $Y2=0
r177 64 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=4.08
+ $Y2=0
r178 63 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r179 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r180 60 63 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r181 60 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r182 59 62 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r183 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r184 57 95 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.747 $Y2=0
r185 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r186 56 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.57
+ $Y2=0
r187 56 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=0
+ $X2=3.12 $Y2=0
r188 54 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r189 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r190 51 95 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.747
+ $Y2=0
r191 51 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.24
+ $Y2=0
r192 49 76 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=8.4
+ $Y2=0
r193 49 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.48 $Y2=0
r194 47 75 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.49 $Y=0 $X2=8.4
+ $Y2=0
r195 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.49 $Y=0 $X2=8.655
+ $Y2=0
r196 46 79 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=8.82 $Y=0 $X2=8.88
+ $Y2=0
r197 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.82 $Y=0 $X2=8.655
+ $Y2=0
r198 44 69 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=6
+ $Y2=0
r199 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=6.31
+ $Y2=0
r200 43 72 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.48
+ $Y2=0
r201 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.31
+ $Y2=0
r202 39 104 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=12.745 $Y=0.085
+ $X2=12.745 $Y2=0
r203 39 41 9.66018 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=12.745 $Y=0.085
+ $X2=12.745 $Y2=0.37
r204 35 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0
r205 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0.38
r206 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.655 $Y=0.085
+ $X2=8.655 $Y2=0
r207 31 33 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=8.655 $Y=0.085
+ $X2=8.655 $Y2=0.8
r208 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.31 $Y=0.085
+ $X2=6.31 $Y2=0
r209 27 29 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=6.31 $Y=0.085
+ $X2=6.31 $Y2=0.775
r210 23 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r211 23 25 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.55
r212 19 95 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0
r213 19 21 17.189 $w=2.93e-07 $l=4.4e-07 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0.525
r214 6 41 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=12.53
+ $Y=0.235 $X2=12.75 $Y2=0.37
r215 5 37 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=10.7
+ $Y=0.785 $X2=10.92 $Y2=0.38
r216 4 33 182 $w=1.7e-07 $l=4.00625e-07 $layer=licon1_NDIFF $count=1 $X=8.355
+ $Y=0.565 $X2=8.655 $Y2=0.8
r217 3 29 182 $w=1.7e-07 $l=4.68375e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.565 $X2=6.31 $Y2=0.775
r218 2 25 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.405 $X2=3.57 $Y2=0.55
r219 1 21 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_OV2%noxref_24 1 2 7 9 14
c28 7 0 1.6277e-19 $X=2.895 $Y=0.35
r29 14 17 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.06 $Y=0.35
+ $X2=3.06 $Y2=0.53
r30 9 12 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.25 $Y=0.35 $X2=1.25
+ $Y2=0.43
r31 8 9 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.355 $Y=0.35 $X2=1.25
+ $Y2=0.35
r32 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0.35
+ $X2=3.06 $Y2=0.35
r33 7 8 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=2.895 $Y=0.35
+ $X2=1.355 $Y2=0.35
r34 2 17 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.92
+ $Y=0.405 $X2=3.06 $Y2=0.53
r35 1 12 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.25 $X2=1.25 $Y2=0.43
.ends

