# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfsbp_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdfsbp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.32000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.460000 2.300000 1.790000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.615000 1.850000 16.210000 2.890000 ;
        RECT 15.880000 0.350000 16.210000 0.810000 ;
        RECT 16.040000 0.810000 16.210000 1.850000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.565000 0.265000 14.075000 0.725000 ;
        RECT 13.565000 0.725000 13.795000 1.610000 ;
        RECT 13.565000 1.610000 14.245000 1.780000 ;
        RECT 13.995000 1.780000 14.245000 3.020000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.110000 3.685000 1.780000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 0.855000 2.275000 1.110000 ;
        RECT 0.930000 1.110000 2.835000 1.185000 ;
        RECT 1.565000 0.810000 2.275000 0.855000 ;
        RECT 1.565000 1.185000 2.835000 1.280000 ;
        RECT 2.510000 1.280000 2.835000 1.790000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  8.735000 1.550000  9.025000 1.595000 ;
        RECT  8.735000 1.595000 12.385000 1.735000 ;
        RECT  8.735000 1.735000  9.025000 1.780000 ;
        RECT 12.095000 1.550000 12.385000 1.595000 ;
        RECT 12.095000 1.735000 12.385000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.215000 1.450000 4.645000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 16.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.320000 0.085000 ;
      RECT  0.000000  3.245000 16.320000 3.415000 ;
      RECT  0.115000  0.265000  0.565000 1.425000 ;
      RECT  0.115000  1.425000  1.385000 1.755000 ;
      RECT  0.115000  1.755000  0.445000 3.065000 ;
      RECT  0.645000  2.025000  0.975000 3.245000 ;
      RECT  1.055000  0.085000  1.385000 0.675000 ;
      RECT  1.205000  2.025000  1.535000 2.895000 ;
      RECT  1.205000  2.895000  2.575000 3.065000 ;
      RECT  1.735000  1.970000  3.185000 2.140000 ;
      RECT  1.735000  2.140000  2.065000 2.715000 ;
      RECT  2.175000  0.265000  2.625000 0.630000 ;
      RECT  2.405000  2.320000  3.615000 2.490000 ;
      RECT  2.405000  2.490000  2.575000 2.895000 ;
      RECT  2.455000  0.630000  2.625000 0.760000 ;
      RECT  2.455000  0.760000  3.675000 0.930000 ;
      RECT  2.755000  2.670000  3.085000 3.245000 ;
      RECT  2.995000  0.085000  3.325000 0.580000 ;
      RECT  3.015000  0.930000  3.185000 1.970000 ;
      RECT  3.285000  2.490000  3.615000 3.065000 ;
      RECT  3.505000  0.265000  4.465000 0.435000 ;
      RECT  3.505000  0.435000  3.675000 0.760000 ;
      RECT  3.850000  1.960000  5.140000 2.130000 ;
      RECT  3.850000  2.130000  4.180000 3.065000 ;
      RECT  3.865000  0.615000  4.115000 1.005000 ;
      RECT  3.865000  1.005000  4.035000 1.960000 ;
      RECT  4.295000  0.435000  4.465000 1.100000 ;
      RECT  4.295000  1.100000  5.185000 1.185000 ;
      RECT  4.295000  1.185000  5.490000 1.270000 ;
      RECT  4.380000  2.310000  4.710000 3.245000 ;
      RECT  4.655000  0.085000  4.825000 0.920000 ;
      RECT  4.825000  1.555000  5.140000 1.960000 ;
      RECT  4.910000  2.310000  5.240000 2.895000 ;
      RECT  4.910000  2.895000  7.560000 3.065000 ;
      RECT  5.015000  0.265000  6.270000 0.435000 ;
      RECT  5.015000  0.435000  5.185000 1.100000 ;
      RECT  5.015000  1.270000  5.490000 1.355000 ;
      RECT  5.320000  1.355000  5.490000 1.960000 ;
      RECT  5.320000  1.960000  5.780000 2.130000 ;
      RECT  5.365000  0.615000  5.840000 1.005000 ;
      RECT  5.450000  2.130000  5.780000 2.715000 ;
      RECT  5.670000  1.005000  5.840000 1.300000 ;
      RECT  5.670000  1.300000  6.905000 1.630000 ;
      RECT  5.670000  1.630000  6.130000 1.780000 ;
      RECT  5.960000  1.780000  6.130000 2.895000 ;
      RECT  6.020000  0.435000  6.270000 0.855000 ;
      RECT  6.310000  2.075000  7.255000 2.245000 ;
      RECT  6.310000  2.245000  6.640000 2.715000 ;
      RECT  6.450000  0.605000  6.780000 0.875000 ;
      RECT  6.450000  0.875000  7.915000 1.045000 ;
      RECT  6.450000  1.045000  6.780000 1.065000 ;
      RECT  7.085000  1.045000  7.255000 2.075000 ;
      RECT  7.315000  0.085000  7.565000 0.695000 ;
      RECT  7.390000  2.515000  9.985000 2.685000 ;
      RECT  7.390000  2.685000  7.560000 2.895000 ;
      RECT  7.435000  1.225000  8.265000 1.395000 ;
      RECT  7.435000  1.395000  7.765000 2.085000 ;
      RECT  7.435000  2.085000  8.600000 2.335000 ;
      RECT  7.740000  2.865000  8.070000 3.245000 ;
      RECT  7.745000  0.265000  8.870000 0.435000 ;
      RECT  7.745000  0.435000  7.915000 0.875000 ;
      RECT  8.005000  1.575000  8.615000 1.905000 ;
      RECT  8.095000  0.615000  8.520000 1.020000 ;
      RECT  8.095000  1.020000  8.265000 1.225000 ;
      RECT  8.445000  1.200000  9.605000 1.370000 ;
      RECT  8.445000  1.370000  8.615000 1.575000 ;
      RECT  8.700000  0.435000  8.870000 1.200000 ;
      RECT  8.795000  1.550000  9.065000 1.880000 ;
      RECT  8.800000  2.865000  9.130000 3.245000 ;
      RECT  9.050000  0.085000  9.380000 1.020000 ;
      RECT  9.275000  1.370000  9.605000 1.870000 ;
      RECT  9.815000  1.155000 10.145000 1.605000 ;
      RECT  9.815000  1.605000 10.980000 1.775000 ;
      RECT  9.815000  1.775000  9.985000 2.515000 ;
      RECT 10.205000  2.075000 10.535000 2.115000 ;
      RECT 10.205000  2.115000 12.460000 2.285000 ;
      RECT 10.205000  2.285000 10.535000 3.065000 ;
      RECT 10.325000  0.310000 10.655000 0.950000 ;
      RECT 10.325000  0.950000 11.330000 1.120000 ;
      RECT 10.715000  1.775000 10.980000 1.935000 ;
      RECT 11.160000  1.120000 11.330000 2.115000 ;
      RECT 11.510000  1.200000 12.810000 1.370000 ;
      RECT 11.510000  1.370000 11.775000 1.885000 ;
      RECT 11.510000  2.465000 11.840000 3.245000 ;
      RECT 11.590000  0.085000 11.920000 0.770000 ;
      RECT 11.985000  1.550000 12.355000 1.890000 ;
      RECT 12.165000  0.265000 12.495000 1.200000 ;
      RECT 12.210000  2.075000 12.460000 2.115000 ;
      RECT 12.210000  2.285000 12.460000 2.895000 ;
      RECT 12.210000  2.895000 13.365000 3.065000 ;
      RECT 12.640000  1.370000 12.810000 2.020000 ;
      RECT 12.640000  2.020000 13.015000 2.715000 ;
      RECT 12.955000  0.085000 13.285000 0.725000 ;
      RECT 12.990000  1.170000 13.365000 1.840000 ;
      RECT 13.195000  1.840000 13.365000 2.895000 ;
      RECT 13.545000  1.980000 13.795000 3.245000 ;
      RECT 14.300000  0.350000 14.630000 0.810000 ;
      RECT 14.460000  0.810000 14.630000 1.490000 ;
      RECT 14.460000  1.490000 15.725000 1.660000 ;
      RECT 14.460000  1.660000 14.885000 2.890000 ;
      RECT 15.085000  1.850000 15.415000 3.245000 ;
      RECT 15.090000  0.085000 15.420000 0.810000 ;
      RECT 15.395000  0.990000 15.725000 1.490000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.580000  8.965000 1.750000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  1.580000 12.325000 1.750000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfsbp_lp
END LIBRARY
