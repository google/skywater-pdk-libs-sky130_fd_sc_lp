* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_1741_137# a_1649_512# VPB phighvt w=420000u l=150000u
+  ad=2.95378e+12p pd=2.258e+07u as=2.709e+11p ps=2.13e+06u
M1001 a_1741_137# a_1531_428# a_1896_119# VNB nshort w=640000u l=150000u
+  ad=2.4475e+11p pd=2.35e+06u as=4.352e+11p ps=3.92e+06u
M1002 VGND RESET_B a_1186_21# VNB nshort w=420000u l=150000u
+  ad=1.9425e+12p pd=1.556e+07u as=1.197e+11p ps=1.41e+06u
M1003 a_1228_379# a_546_449# a_755_398# VPB phighvt w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=7.14e+11p ps=3.38e+06u
M1004 a_1436_379# a_755_398# VPWR VPB phighvt w=840000u l=150000u
+  ad=3.15875e+11p pd=2.82e+06u as=0p ps=0u
M1005 a_1442_119# a_755_398# VGND VNB nshort w=640000u l=150000u
+  ad=2.304e+11p pd=2e+06u as=0p ps=0u
M1006 VGND a_1741_137# a_1693_163# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 VPWR RESET_B a_1186_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1008 a_460_449# D VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1009 VGND a_113_67# a_223_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1010 VPWR a_755_398# a_707_449# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1011 Q_N a_1741_137# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.465e+11p pd=3.07e+06u as=0p ps=0u
M1012 a_1013_66# a_1186_21# a_755_398# VNB nshort w=640000u l=150000u
+  ad=3.648e+11p pd=3.7e+06u as=3.606e+11p ps=2.75e+06u
M1013 VPWR a_1186_21# a_2036_451# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1014 a_1896_119# a_1186_21# a_1741_137# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1741_137# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 Q a_2511_137# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1017 a_755_398# a_546_449# a_1013_66# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1693_163# a_223_119# a_1531_428# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.643e+11p ps=2.47e+06u
M1019 VPWR a_1741_137# a_2511_137# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1020 VPWR a_1186_21# a_1228_379# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1531_428# a_223_119# a_1436_379# VPB phighvt w=840000u l=150000u
+  ad=3.381e+11p pd=2.56e+06u as=0p ps=0u
M1022 a_460_449# D VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1023 a_546_449# a_223_119# a_460_449# VNB nshort w=420000u l=150000u
+  ad=2.2095e+11p pd=1.92e+06u as=0p ps=0u
M1024 a_1013_66# SET_B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1531_428# a_113_67# a_1442_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1896_119# SET_B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_113_67# CLK_N VPWR VPB phighvt w=640000u l=150000u
+  ad=2.336e+11p pd=2.01e+06u as=0p ps=0u
M1028 a_2036_451# a_1531_428# a_1741_137# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_113_67# CLK_N VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1030 Q_N a_1741_137# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1031 VGND a_755_398# a_702_110# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1032 VPWR a_113_67# a_223_119# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1033 a_707_449# a_223_119# a_546_449# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.751e+11p ps=2.15e+06u
M1034 VGND a_1741_137# a_2511_137# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1035 Q a_2511_137# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1036 a_546_449# a_113_67# a_460_449# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_755_398# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_702_110# a_113_67# a_546_449# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1649_512# a_113_67# a_1531_428# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
