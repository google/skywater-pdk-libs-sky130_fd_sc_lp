* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VGND A3 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_192_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND A2 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_192_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_981_361# A3 a_554_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A1 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_554_361# A3 a_981_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_1346_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND A3 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_1346_367# A2 a_981_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_192_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_554_361# A3 a_981_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_192_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR A1 a_1346_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_192_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Y B1 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_192_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_981_361# A2 a_1346_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_192_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 VGND A2 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_192_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Y B1 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_981_361# A2 a_1346_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_554_361# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_1346_367# A2 a_981_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_192_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 Y A4 a_554_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VGND A4 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 VGND A4 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_192_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 a_981_361# A3 a_554_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 VPWR A1 a_1346_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 VGND A1 a_192_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 Y A4 a_554_361# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 a_1346_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 a_554_361# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
