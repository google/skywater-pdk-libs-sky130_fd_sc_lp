* File: sky130_fd_sc_lp__o2111a_0.pxi.spice
* Created: Wed Sep  2 10:12:08 2020
* 
x_PM_SKY130_FD_SC_LP__O2111A_0%A_80_21# N_A_80_21#_M1001_s N_A_80_21#_M1008_d
+ N_A_80_21#_M1011_d N_A_80_21#_M1003_g N_A_80_21#_c_95_n N_A_80_21#_M1002_g
+ N_A_80_21#_c_97_n N_A_80_21#_c_90_n N_A_80_21#_c_91_n N_A_80_21#_c_92_n
+ N_A_80_21#_c_93_n N_A_80_21#_c_99_n N_A_80_21#_c_100_n N_A_80_21#_c_94_n
+ N_A_80_21#_c_101_n N_A_80_21#_c_102_n N_A_80_21#_c_103_n N_A_80_21#_c_104_n
+ PM_SKY130_FD_SC_LP__O2111A_0%A_80_21#
x_PM_SKY130_FD_SC_LP__O2111A_0%D1 N_D1_M1008_g N_D1_c_180_n N_D1_M1001_g
+ N_D1_c_181_n N_D1_c_182_n N_D1_c_183_n N_D1_c_184_n D1 D1 N_D1_c_186_n
+ PM_SKY130_FD_SC_LP__O2111A_0%D1
x_PM_SKY130_FD_SC_LP__O2111A_0%C1 N_C1_c_235_n N_C1_M1000_g N_C1_M1004_g
+ N_C1_c_237_n C1 C1 C1 C1 N_C1_c_239_n PM_SKY130_FD_SC_LP__O2111A_0%C1
x_PM_SKY130_FD_SC_LP__O2111A_0%B1 N_B1_M1005_g N_B1_c_285_n N_B1_M1011_g
+ N_B1_c_290_n B1 B1 N_B1_c_287_n PM_SKY130_FD_SC_LP__O2111A_0%B1
x_PM_SKY130_FD_SC_LP__O2111A_0%A2 N_A2_c_325_n N_A2_M1010_g N_A2_M1006_g
+ N_A2_c_326_n N_A2_c_327_n N_A2_c_328_n N_A2_c_332_n A2 A2 N_A2_c_330_n
+ PM_SKY130_FD_SC_LP__O2111A_0%A2
x_PM_SKY130_FD_SC_LP__O2111A_0%A1 N_A1_c_375_n N_A1_M1009_g N_A1_M1007_g
+ N_A1_c_376_n N_A1_c_377_n N_A1_c_378_n N_A1_c_383_n N_A1_c_379_n A1 A1 A1
+ N_A1_c_380_n PM_SKY130_FD_SC_LP__O2111A_0%A1
x_PM_SKY130_FD_SC_LP__O2111A_0%X N_X_M1003_s N_X_M1002_s X X X X X X X
+ N_X_c_415_n X PM_SKY130_FD_SC_LP__O2111A_0%X
x_PM_SKY130_FD_SC_LP__O2111A_0%VPWR N_VPWR_M1002_d N_VPWR_M1000_d N_VPWR_M1007_d
+ N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n
+ N_VPWR_c_438_n VPWR N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n
+ N_VPWR_c_432_n PM_SKY130_FD_SC_LP__O2111A_0%VPWR
x_PM_SKY130_FD_SC_LP__O2111A_0%VGND N_VGND_M1003_d N_VGND_M1010_d N_VGND_c_476_n
+ N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n VGND N_VGND_c_480_n
+ N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n PM_SKY130_FD_SC_LP__O2111A_0%VGND
x_PM_SKY130_FD_SC_LP__O2111A_0%A_459_47# N_A_459_47#_M1005_d N_A_459_47#_M1009_d
+ N_A_459_47#_c_533_n N_A_459_47#_c_534_n N_A_459_47#_c_535_n
+ N_A_459_47#_c_536_n PM_SKY130_FD_SC_LP__O2111A_0%A_459_47#
cc_1 VNB N_A_80_21#_M1003_g 0.0678884f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_80_21#_c_90_n 0.00646611f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.71
cc_3 VNB N_A_80_21#_c_91_n 0.0161269f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.71
cc_4 VNB N_A_80_21#_c_92_n 0.0152133f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.825
cc_5 VNB N_A_80_21#_c_93_n 0.00254042f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=0.825
cc_6 VNB N_A_80_21#_c_94_n 0.00615905f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.445
cc_7 VNB N_D1_c_180_n 0.0181234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D1_c_181_n 0.0113201f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_9 VNB N_D1_c_182_n 0.0259111f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_10 VNB N_D1_c_183_n 0.00486169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_D1_c_184_n 0.0272476f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.215
cc_12 VNB D1 0.00167913f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.725
cc_13 VNB N_D1_c_186_n 0.0184712f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.71
cc_14 VNB N_C1_c_235_n 0.0200061f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=2.405
cc_15 VNB N_C1_M1004_g 0.033061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_c_237_n 6.49549e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_17 VNB C1 0.00531428f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_18 VNB N_C1_c_239_n 0.0176853f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.91
cc_19 VNB N_B1_M1005_g 0.0375363f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.405
cc_20 VNB N_B1_c_285_n 0.0163357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB B1 0.0137115f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_22 VNB N_B1_c_287_n 0.0165326f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.725
cc_23 VNB N_A2_c_325_n 0.0164575f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.235
cc_24 VNB N_A2_c_326_n 0.020496f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_25 VNB N_A2_c_327_n 0.0153602f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=2.018
cc_26 VNB N_A2_c_328_n 0.0215546f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.215
cc_27 VNB A2 0.00646808f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.725
cc_28 VNB N_A2_c_330_n 0.0160848f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.71
cc_29 VNB N_A1_c_375_n 0.0201853f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.235
cc_30 VNB N_A1_c_376_n 0.0654536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A1_c_377_n 0.0241303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_c_378_n 0.00182823f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_33 VNB N_A1_c_379_n 0.0251435f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.215
cc_34 VNB N_A1_c_380_n 0.0250208f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.825
cc_35 VNB N_X_c_415_n 0.0673492f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.71
cc_36 VNB N_VPWR_c_432_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.71
cc_37 VNB N_VGND_c_476_n 0.00686958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_477_n 0.00561441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_478_n 0.0509231f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.215
cc_40 VNB N_VGND_c_479_n 0.00631792f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.725
cc_41 VNB N_VGND_c_480_n 0.0153306f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=2.215
cc_42 VNB N_VGND_c_481_n 0.0235765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_482_n 0.22082f $X=-0.19 $Y=-0.245 $X2=1.437 $Y2=2.215
cc_44 VNB N_VGND_c_483_n 0.00510715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_459_47#_c_533_n 3.66741e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_459_47#_c_534_n 0.0127778f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_47 VNB N_A_459_47#_c_535_n 0.00384408f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_48 VNB N_A_459_47#_c_536_n 0.0162223f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=2.018
cc_49 VPB N_A_80_21#_c_95_n 0.0239644f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=2.018
cc_50 VPB N_A_80_21#_M1002_g 0.0257408f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.725
cc_51 VPB N_A_80_21#_c_97_n 0.0228216f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=2.215
cc_52 VPB N_A_80_21#_c_91_n 0.00724709f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.71
cc_53 VPB N_A_80_21#_c_99_n 0.0139927f $X=-0.19 $Y=1.655 $X2=1.305 $Y2=2.125
cc_54 VPB N_A_80_21#_c_100_n 0.00112463f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.125
cc_55 VPB N_A_80_21#_c_101_n 0.0060826f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=2.55
cc_56 VPB N_A_80_21#_c_102_n 0.0242593f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=2.125
cc_57 VPB N_A_80_21#_c_103_n 0.00395345f $X=-0.19 $Y=1.655 $X2=2.635 $Y2=2.55
cc_58 VPB N_A_80_21#_c_104_n 0.00802257f $X=-0.19 $Y=1.655 $X2=1.437 $Y2=2.125
cc_59 VPB N_D1_M1008_g 0.0451326f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=2.405
cc_60 VPB N_D1_c_183_n 0.0117052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB D1 0.00316491f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.725
cc_62 VPB N_C1_M1000_g 0.0468308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_C1_c_237_n 0.0171332f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_64 VPB C1 0.00308176f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_65 VPB N_B1_c_285_n 0.00169797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_B1_M1011_g 0.044916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_B1_c_290_n 0.0169607f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_68 VPB B1 0.00595256f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_69 VPB N_A2_M1006_g 0.0397815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A2_c_332_n 0.0157573f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.725
cc_71 VPB A2 0.011118f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.725
cc_72 VPB N_A1_M1007_g 0.0269148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A1_c_378_n 0.0268823f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_74 VPB N_A1_c_383_n 0.0244675f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.742
cc_75 VPB N_A1_c_380_n 0.0301069f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=0.825
cc_76 VPB N_X_c_415_n 0.0386506f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.71
cc_77 VPB X 0.0427802f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=2.125
cc_78 VPB N_VPWR_c_433_n 0.00901792f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_79 VPB N_VPWR_c_434_n 0.013799f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.215
cc_80 VPB N_VPWR_c_435_n 0.0156631f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.725
cc_81 VPB N_VPWR_c_436_n 0.0337924f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=2.215
cc_82 VPB N_VPWR_c_437_n 0.0234952f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.71
cc_83 VPB N_VPWR_c_438_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.71
cc_84 VPB N_VPWR_c_439_n 0.0167145f $X=-0.19 $Y=1.655 $X2=1.247 $Y2=0.445
cc_85 VPB N_VPWR_c_440_n 0.0255809f $X=-0.19 $Y=1.655 $X2=1.437 $Y2=2.55
cc_86 VPB N_VPWR_c_441_n 0.011515f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=2.55
cc_87 VPB N_VPWR_c_432_n 0.0707955f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.71
cc_88 N_A_80_21#_c_95_n N_D1_M1008_g 0.0275486f $X=0.597 $Y=2.018 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_90_n N_D1_M1008_g 0.00113401f $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_99_n N_D1_M1008_g 0.0158f $X=1.305 $Y=2.125 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_101_n N_D1_M1008_g 0.00504726f $X=1.435 $Y=2.55 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_92_n N_D1_c_180_n 5.60297e-19 $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_94_n N_D1_c_180_n 0.00218198f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_90_n N_D1_c_182_n 7.51687e-19 $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_91_n N_D1_c_182_n 0.00535295f $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_95_n N_D1_c_183_n 0.00535295f $X=0.597 $Y=2.018 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_99_n N_D1_c_183_n 6.19693e-19 $X=1.305 $Y=2.125 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_104_n N_D1_c_183_n 5.74242e-19 $X=1.437 $Y=2.125 $X2=0 $Y2=0
cc_99 N_A_80_21#_M1003_g N_D1_c_184_n 0.00345888f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_90_n N_D1_c_184_n 0.00325594f $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_92_n N_D1_c_184_n 0.0134551f $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_102 N_A_80_21#_M1003_g D1 4.27272e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_95_n D1 8.60918e-19 $X=0.597 $Y=2.018 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_90_n D1 0.0463052f $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_91_n D1 7.77022e-19 $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_92_n D1 0.0272139f $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_99_n D1 0.0215226f $X=1.305 $Y=2.125 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_104_n D1 0.00505924f $X=1.437 $Y=2.125 $X2=0 $Y2=0
cc_109 N_A_80_21#_M1003_g N_D1_c_186_n 0.00900676f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_90_n N_D1_c_186_n 0.0039713f $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_92_n N_D1_c_186_n 0.00131738f $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_101_n N_C1_M1000_g 0.00508139f $X=1.435 $Y=2.55 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_102_n N_C1_M1000_g 0.0168127f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_102_n N_C1_c_237_n 0.00404455f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_92_n C1 0.0135842f $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_94_n C1 0.0168862f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_102_n C1 0.0227936f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_104_n C1 0.00224874f $X=1.437 $Y=2.125 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_102_n N_B1_M1011_g 0.0168127f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_103_n N_B1_M1011_g 0.00509728f $X=2.635 $Y=2.55 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_102_n N_B1_c_290_n 0.00146722f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_102_n B1 0.0387523f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_102_n N_A2_M1006_g 0.00579617f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_103_n N_A2_M1006_g 0.0161914f $X=2.635 $Y=2.55 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_102_n N_A2_c_332_n 4.49908e-19 $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_102_n A2 0.00627038f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_103_n N_A1_M1007_g 0.00272933f $X=2.635 $Y=2.55 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_102_n N_A1_c_383_n 5.20657e-19 $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_102_n N_A1_c_380_n 0.00475737f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_130 N_A_80_21#_M1003_g N_X_c_415_n 0.0401512f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_80_21#_M1002_g N_X_c_415_n 0.00537893f $X=0.72 $Y=2.725 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_90_n N_X_c_415_n 0.0861582f $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_133 N_A_80_21#_c_93_n N_X_c_415_n 0.0140511f $X=0.795 $Y=0.825 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_100_n N_X_c_415_n 0.0148776f $X=0.795 $Y=2.125 $X2=0 $Y2=0
cc_135 N_A_80_21#_M1002_g X 0.00836093f $X=0.72 $Y=2.725 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_97_n X 0.00694355f $X=0.597 $Y=2.215 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_100_n X 0.0127302f $X=0.795 $Y=2.125 $X2=0 $Y2=0
cc_138 N_A_80_21#_M1002_g N_VPWR_c_433_n 0.00293165f $X=0.72 $Y=2.725 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_c_99_n N_VPWR_c_433_n 0.0248436f $X=1.305 $Y=2.125 $X2=0 $Y2=0
cc_140 N_A_80_21#_c_101_n N_VPWR_c_433_n 0.00389517f $X=1.435 $Y=2.55 $X2=0
+ $Y2=0
cc_141 N_A_80_21#_c_101_n N_VPWR_c_434_n 0.00411749f $X=1.435 $Y=2.55 $X2=0
+ $Y2=0
cc_142 N_A_80_21#_c_102_n N_VPWR_c_434_n 0.0507046f $X=2.51 $Y=2.125 $X2=0 $Y2=0
cc_143 N_A_80_21#_c_103_n N_VPWR_c_434_n 0.00414404f $X=2.635 $Y=2.55 $X2=0
+ $Y2=0
cc_144 N_A_80_21#_c_103_n N_VPWR_c_436_n 0.0228594f $X=2.635 $Y=2.55 $X2=0 $Y2=0
cc_145 N_A_80_21#_M1002_g N_VPWR_c_437_n 0.00502664f $X=0.72 $Y=2.725 $X2=0
+ $Y2=0
cc_146 N_A_80_21#_c_101_n N_VPWR_c_439_n 0.0188536f $X=1.435 $Y=2.55 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_103_n N_VPWR_c_440_n 0.0205614f $X=2.635 $Y=2.55 $X2=0 $Y2=0
cc_148 N_A_80_21#_M1002_g N_VPWR_c_432_n 0.0102782f $X=0.72 $Y=2.725 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_101_n N_VPWR_c_432_n 0.0102248f $X=1.435 $Y=2.55 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_103_n N_VPWR_c_432_n 0.011087f $X=2.635 $Y=2.55 $X2=0 $Y2=0
cc_151 N_A_80_21#_M1003_g N_VGND_c_476_n 0.0108284f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_152 N_A_80_21#_c_92_n N_VGND_c_476_n 0.00473912f $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_93_n N_VGND_c_476_n 0.0210138f $X=0.795 $Y=0.825 $X2=0 $Y2=0
cc_154 N_A_80_21#_c_94_n N_VGND_c_476_n 0.0173938f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A_80_21#_c_92_n N_VGND_c_478_n 0.00390094f $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_156 N_A_80_21#_c_94_n N_VGND_c_478_n 0.015111f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A_80_21#_M1003_g N_VGND_c_480_n 0.00486043f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_158 N_A_80_21#_M1001_s N_VGND_c_482_n 0.00276582f $X=1.16 $Y=0.235 $X2=0
+ $Y2=0
cc_159 N_A_80_21#_M1003_g N_VGND_c_482_n 0.0093594f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_160 N_A_80_21#_c_92_n N_VGND_c_482_n 0.00723096f $X=1.12 $Y=0.825 $X2=0 $Y2=0
cc_161 N_A_80_21#_c_93_n N_VGND_c_482_n 0.00113336f $X=0.795 $Y=0.825 $X2=0
+ $Y2=0
cc_162 N_A_80_21#_c_94_n N_VGND_c_482_n 0.00969541f $X=1.285 $Y=0.445 $X2=0
+ $Y2=0
cc_163 N_D1_c_182_n N_C1_c_235_n 0.0123814f $X=1.2 $Y=1.585 $X2=0 $Y2=0
cc_164 N_D1_c_180_n N_C1_M1004_g 0.0524924f $X=1.5 $Y=0.765 $X2=0 $Y2=0
cc_165 N_D1_c_181_n N_C1_M1004_g 0.00553277f $X=1.2 $Y=1.08 $X2=0 $Y2=0
cc_166 N_D1_M1008_g N_C1_c_237_n 0.0344949f $X=1.22 $Y=2.725 $X2=0 $Y2=0
cc_167 N_D1_c_183_n N_C1_c_237_n 0.0123814f $X=1.2 $Y=1.75 $X2=0 $Y2=0
cc_168 D1 N_C1_c_237_n 3.81882e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_169 N_D1_M1008_g C1 3.50385e-19 $X=1.22 $Y=2.725 $X2=0 $Y2=0
cc_170 N_D1_c_180_n C1 0.00819572f $X=1.5 $Y=0.765 $X2=0 $Y2=0
cc_171 N_D1_c_181_n C1 0.00800796f $X=1.2 $Y=1.08 $X2=0 $Y2=0
cc_172 N_D1_c_184_n C1 0.00474788f $X=1.5 $Y=0.84 $X2=0 $Y2=0
cc_173 D1 C1 0.0583573f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_174 D1 N_C1_c_239_n 6.95286e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_175 N_D1_c_186_n N_C1_c_239_n 0.0123814f $X=1.2 $Y=1.245 $X2=0 $Y2=0
cc_176 N_D1_M1008_g N_VPWR_c_433_n 0.00180461f $X=1.22 $Y=2.725 $X2=0 $Y2=0
cc_177 N_D1_M1008_g N_VPWR_c_439_n 0.0053602f $X=1.22 $Y=2.725 $X2=0 $Y2=0
cc_178 N_D1_M1008_g N_VPWR_c_432_n 0.0103302f $X=1.22 $Y=2.725 $X2=0 $Y2=0
cc_179 N_D1_c_180_n N_VGND_c_476_n 0.00301907f $X=1.5 $Y=0.765 $X2=0 $Y2=0
cc_180 N_D1_c_180_n N_VGND_c_478_n 0.00545968f $X=1.5 $Y=0.765 $X2=0 $Y2=0
cc_181 N_D1_c_184_n N_VGND_c_478_n 0.00113713f $X=1.5 $Y=0.84 $X2=0 $Y2=0
cc_182 N_D1_c_180_n N_VGND_c_482_n 0.0111542f $X=1.5 $Y=0.765 $X2=0 $Y2=0
cc_183 N_D1_c_184_n N_VGND_c_482_n 0.001077f $X=1.5 $Y=0.84 $X2=0 $Y2=0
cc_184 N_C1_M1004_g N_B1_M1005_g 0.0261227f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_185 C1 N_B1_M1005_g 0.00354875f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_186 N_C1_c_235_n N_B1_c_285_n 0.0261227f $X=1.755 $Y=1.645 $X2=0 $Y2=0
cc_187 N_C1_M1000_g N_B1_M1011_g 0.0128355f $X=1.65 $Y=2.725 $X2=0 $Y2=0
cc_188 N_C1_M1000_g N_B1_c_290_n 0.00101856f $X=1.65 $Y=2.725 $X2=0 $Y2=0
cc_189 N_C1_c_237_n N_B1_c_290_n 0.0261227f $X=1.755 $Y=1.825 $X2=0 $Y2=0
cc_190 N_C1_M1004_g B1 0.00475888f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_191 C1 B1 0.0589703f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_192 N_C1_c_239_n N_B1_c_287_n 0.0261227f $X=1.77 $Y=1.32 $X2=0 $Y2=0
cc_193 N_C1_M1000_g N_VPWR_c_434_n 0.00234444f $X=1.65 $Y=2.725 $X2=0 $Y2=0
cc_194 N_C1_M1000_g N_VPWR_c_439_n 0.0053602f $X=1.65 $Y=2.725 $X2=0 $Y2=0
cc_195 N_C1_M1000_g N_VPWR_c_432_n 0.0106597f $X=1.65 $Y=2.725 $X2=0 $Y2=0
cc_196 N_C1_M1004_g N_VGND_c_478_n 0.00491601f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_197 C1 N_VGND_c_478_n 0.00986007f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_198 N_C1_M1004_g N_VGND_c_482_n 0.00812684f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_199 C1 N_VGND_c_482_n 0.0107248f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_200 C1 A_315_47# 0.00119247f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_201 N_C1_M1004_g N_A_459_47#_c_533_n 0.00132552f $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_202 C1 N_A_459_47#_c_533_n 0.0115109f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_203 N_C1_M1004_g N_A_459_47#_c_535_n 4.48779e-19 $X=1.86 $Y=0.445 $X2=0 $Y2=0
cc_204 C1 N_A_459_47#_c_535_n 0.00655497f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_205 N_B1_M1005_g N_A2_c_325_n 0.0198f $X=2.22 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_206 N_B1_M1011_g N_A2_M1006_g 0.0304918f $X=2.42 $Y=2.725 $X2=0 $Y2=0
cc_207 N_B1_c_290_n N_A2_M1006_g 0.00172456f $X=2.325 $Y=1.865 $X2=0 $Y2=0
cc_208 B1 N_A2_M1006_g 9.02196e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_209 N_B1_M1005_g N_A2_c_327_n 0.00918703f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_210 B1 N_A2_c_327_n 0.00420058f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_211 N_B1_c_285_n N_A2_c_328_n 0.013165f $X=2.325 $Y=1.685 $X2=0 $Y2=0
cc_212 N_B1_c_290_n N_A2_c_332_n 0.013165f $X=2.325 $Y=1.865 $X2=0 $Y2=0
cc_213 B1 A2 0.0499703f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_214 N_B1_c_287_n A2 7.81337e-19 $X=2.34 $Y=1.36 $X2=0 $Y2=0
cc_215 N_B1_c_287_n N_A2_c_330_n 0.013165f $X=2.34 $Y=1.36 $X2=0 $Y2=0
cc_216 N_B1_M1011_g N_VPWR_c_434_n 0.00364512f $X=2.42 $Y=2.725 $X2=0 $Y2=0
cc_217 N_B1_M1011_g N_VPWR_c_440_n 0.0053602f $X=2.42 $Y=2.725 $X2=0 $Y2=0
cc_218 N_B1_M1011_g N_VPWR_c_432_n 0.0106324f $X=2.42 $Y=2.725 $X2=0 $Y2=0
cc_219 N_B1_M1005_g N_VGND_c_478_n 0.0054978f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_220 N_B1_M1005_g N_VGND_c_482_n 0.00995168f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_221 N_B1_M1005_g N_A_459_47#_c_533_n 0.00720629f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_222 N_B1_M1005_g N_A_459_47#_c_535_n 0.00502442f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_223 B1 N_A_459_47#_c_535_n 0.0155643f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_224 N_B1_c_287_n N_A_459_47#_c_535_n 0.00135222f $X=2.34 $Y=1.36 $X2=0 $Y2=0
cc_225 N_A2_c_325_n N_A1_c_375_n 0.0102757f $X=2.65 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A2_c_326_n N_A1_c_376_n 0.0102264f $X=2.79 $Y=0.84 $X2=0 $Y2=0
cc_227 N_A2_c_327_n N_A1_c_376_n 0.00765177f $X=2.88 $Y=1.155 $X2=0 $Y2=0
cc_228 A2 N_A1_c_376_n 0.00899606f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_229 N_A2_c_330_n N_A1_c_377_n 0.00988425f $X=2.88 $Y=1.32 $X2=0 $Y2=0
cc_230 N_A2_M1006_g N_A1_c_378_n 0.00751258f $X=2.85 $Y=2.725 $X2=0 $Y2=0
cc_231 N_A2_c_332_n N_A1_c_378_n 0.00988425f $X=2.88 $Y=1.825 $X2=0 $Y2=0
cc_232 N_A2_M1006_g N_A1_c_383_n 0.0655594f $X=2.85 $Y=2.725 $X2=0 $Y2=0
cc_233 A2 N_A1_c_383_n 0.00352551f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_234 N_A2_c_328_n N_A1_c_379_n 0.00988425f $X=2.88 $Y=1.66 $X2=0 $Y2=0
cc_235 N_A2_M1006_g N_A1_c_380_n 0.00146902f $X=2.85 $Y=2.725 $X2=0 $Y2=0
cc_236 N_A2_c_327_n N_A1_c_380_n 5.26092e-19 $X=2.88 $Y=1.155 $X2=0 $Y2=0
cc_237 A2 N_A1_c_380_n 0.0563917f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_238 N_A2_c_330_n N_A1_c_380_n 5.71008e-19 $X=2.88 $Y=1.32 $X2=0 $Y2=0
cc_239 N_A2_M1006_g N_VPWR_c_436_n 0.00268787f $X=2.85 $Y=2.725 $X2=0 $Y2=0
cc_240 N_A2_M1006_g N_VPWR_c_440_n 0.00502372f $X=2.85 $Y=2.725 $X2=0 $Y2=0
cc_241 N_A2_M1006_g N_VPWR_c_432_n 0.00944803f $X=2.85 $Y=2.725 $X2=0 $Y2=0
cc_242 N_A2_c_325_n N_VGND_c_477_n 0.00328698f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_243 N_A2_c_326_n N_VGND_c_477_n 7.12182e-19 $X=2.79 $Y=0.84 $X2=0 $Y2=0
cc_244 N_A2_c_325_n N_VGND_c_478_n 0.00433717f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_245 N_A2_c_325_n N_VGND_c_482_n 0.00606522f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_246 N_A2_c_325_n N_A_459_47#_c_533_n 0.00114558f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_247 N_A2_c_325_n N_A_459_47#_c_534_n 0.00638177f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_248 N_A2_c_326_n N_A_459_47#_c_534_n 0.0147559f $X=2.79 $Y=0.84 $X2=0 $Y2=0
cc_249 A2 N_A_459_47#_c_534_n 0.0282529f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_250 N_A2_c_330_n N_A_459_47#_c_534_n 0.00109866f $X=2.88 $Y=1.32 $X2=0 $Y2=0
cc_251 N_A1_M1007_g N_VPWR_c_436_n 0.0176808f $X=3.21 $Y=2.725 $X2=0 $Y2=0
cc_252 N_A1_c_383_n N_VPWR_c_436_n 0.00683887f $X=3.39 $Y=2.14 $X2=0 $Y2=0
cc_253 N_A1_c_380_n N_VPWR_c_436_n 0.0175439f $X=3.55 $Y=1.12 $X2=0 $Y2=0
cc_254 N_A1_M1007_g N_VPWR_c_440_n 0.00445056f $X=3.21 $Y=2.725 $X2=0 $Y2=0
cc_255 N_A1_M1007_g N_VPWR_c_432_n 0.0079903f $X=3.21 $Y=2.725 $X2=0 $Y2=0
cc_256 N_A1_c_375_n N_VGND_c_477_n 0.00328698f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_257 N_A1_c_375_n N_VGND_c_481_n 0.00433717f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_258 N_A1_c_376_n N_VGND_c_481_n 5.74712e-19 $X=3.515 $Y=1.155 $X2=0 $Y2=0
cc_259 N_A1_c_375_n N_VGND_c_482_n 0.0072035f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_260 N_A1_c_375_n N_A_459_47#_c_534_n 0.00696225f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_261 N_A1_c_376_n N_A_459_47#_c_534_n 0.0232306f $X=3.515 $Y=1.155 $X2=0 $Y2=0
cc_262 N_A1_c_380_n N_A_459_47#_c_534_n 0.0123391f $X=3.55 $Y=1.12 $X2=0 $Y2=0
cc_263 N_A1_c_375_n N_A_459_47#_c_536_n 0.00195506f $X=3.15 $Y=0.765 $X2=0 $Y2=0
cc_264 X N_VPWR_c_433_n 0.0294035f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_265 X N_VPWR_c_437_n 0.0392254f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_266 X N_VPWR_c_432_n 0.0224476f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_267 N_X_c_415_n N_VGND_c_480_n 0.0174138f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_268 N_X_M1003_s N_VGND_c_482_n 0.0037619f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_269 N_X_c_415_n N_VGND_c_482_n 0.0103698f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_270 N_VGND_c_482_n A_315_47# 0.00179454f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_271 N_VGND_c_482_n A_387_47# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_272 N_VGND_c_482_n N_A_459_47#_M1005_d 0.00229771f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_273 N_VGND_c_482_n N_A_459_47#_M1009_d 0.00227158f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_274 N_VGND_c_478_n N_A_459_47#_c_533_n 0.0144931f $X=2.735 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_482_n N_A_459_47#_c_533_n 0.0110829f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_477_n N_A_459_47#_c_534_n 0.0217901f $X=2.9 $Y=0.41 $X2=0 $Y2=0
cc_277 N_VGND_c_478_n N_A_459_47#_c_534_n 0.00244542f $X=2.735 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_481_n N_A_459_47#_c_534_n 0.00268725f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_482_n N_A_459_47#_c_534_n 0.00940437f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_481_n N_A_459_47#_c_536_n 0.0158049f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_c_482_n N_A_459_47#_c_536_n 0.0106312f $X=3.6 $Y=0 $X2=0 $Y2=0
