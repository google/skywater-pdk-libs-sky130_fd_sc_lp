* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a22o_m A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_85_317# B1 a_265_501# VPB phighvt w=420000u l=150000u
+  ad=2.258e+11p pd=1.94e+06u as=2.352e+11p ps=2.8e+06u
M1001 VGND a_85_317# X VNB nshort w=420000u l=150000u
+  ad=3.402e+11p pd=3.3e+06u as=1.197e+11p ps=1.41e+06u
M1002 VPWR a_85_317# X VPB phighvt w=420000u l=150000u
+  ad=3.045e+11p pd=3.13e+06u as=1.113e+11p ps=1.37e+06u
M1003 VPWR A1 a_265_501# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_85_317# A1 a_265_125# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_265_501# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_265_501# B2 a_85_317# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_265_125# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B2 a_445_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 a_445_125# B1 a_85_317# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
