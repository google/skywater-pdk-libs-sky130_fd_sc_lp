# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ha_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__ha_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.495000 0.815000 1.805000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.495000 1.315000 1.795000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 0.255000 3.725000 1.015000 ;
        RECT 3.450000 1.015000 3.725000 2.305000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 1.695000 4.645000 3.075000 ;
        RECT 4.465000 0.255000 4.645000 1.695000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.185000  0.650000 0.515000 1.075000 ;
      RECT 0.185000  1.075000 1.315000 1.245000 ;
      RECT 0.320000  1.975000 0.650000 3.245000 ;
      RECT 0.685000  0.085000 0.935000 0.905000 ;
      RECT 1.105000  0.650000 1.315000 1.075000 ;
      RECT 1.110000  1.965000 1.655000 2.135000 ;
      RECT 1.110000  2.135000 1.390000 2.635000 ;
      RECT 1.485000  0.650000 1.805000 0.980000 ;
      RECT 1.485000  0.980000 1.660000 1.685000 ;
      RECT 1.485000  1.685000 2.335000 1.855000 ;
      RECT 1.485000  1.855000 1.655000 1.965000 ;
      RECT 1.780000  2.255000 1.995000 3.245000 ;
      RECT 1.840000  1.150000 2.335000 1.185000 ;
      RECT 1.840000  1.185000 3.280000 1.515000 ;
      RECT 1.975000  0.700000 2.335000 1.150000 ;
      RECT 2.165000  1.855000 2.335000 2.475000 ;
      RECT 2.165000  2.475000 4.140000 2.645000 ;
      RECT 2.505000  1.515000 2.695000 2.305000 ;
      RECT 2.795000  0.085000 3.220000 1.015000 ;
      RECT 2.950000  2.815000 3.280000 3.245000 ;
      RECT 3.810000  2.815000 4.140000 3.245000 ;
      RECT 3.895000  0.085000 4.225000 1.015000 ;
      RECT 3.970000  1.185000 4.295000 1.515000 ;
      RECT 3.970000  1.515000 4.140000 2.475000 ;
      RECT 4.815000  1.815000 5.015000 3.245000 ;
      RECT 4.825000  0.085000 5.155000 1.095000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_lp__ha_2
END LIBRARY
