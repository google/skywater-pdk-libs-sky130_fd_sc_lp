* File: sky130_fd_sc_lp__xor2_2.pxi.spice
* Created: Fri Aug 28 11:36:21 2020
* 
x_PM_SKY130_FD_SC_LP__XOR2_2%A N_A_M1003_g N_A_M1001_g N_A_M1015_g N_A_M1004_g
+ N_A_M1006_g N_A_M1008_g N_A_M1013_g N_A_M1010_g N_A_c_106_n N_A_c_130_p
+ N_A_c_293_p N_A_c_107_n N_A_c_108_n N_A_c_109_n N_A_c_145_p N_A_c_202_p
+ N_A_c_125_n N_A_c_110_n N_A_c_111_n N_A_c_236_p N_A_c_112_n N_A_c_113_n A A
+ N_A_c_114_n N_A_c_115_n N_A_c_116_n N_A_c_117_n N_A_c_118_n
+ PM_SKY130_FD_SC_LP__XOR2_2%A
x_PM_SKY130_FD_SC_LP__XOR2_2%B N_B_M1009_g N_B_M1000_g N_B_M1014_g N_B_M1011_g
+ N_B_M1012_g N_B_M1005_g N_B_M1018_g N_B_M1017_g N_B_c_328_n N_B_c_337_n B
+ N_B_c_329_n N_B_c_330_n N_B_c_341_n N_B_c_331_n PM_SKY130_FD_SC_LP__XOR2_2%B
x_PM_SKY130_FD_SC_LP__XOR2_2%A_149_65# N_A_149_65#_M1003_s N_A_149_65#_M1011_s
+ N_A_149_65#_M1000_s N_A_149_65#_c_467_n N_A_149_65#_M1007_g
+ N_A_149_65#_M1002_g N_A_149_65#_c_469_n N_A_149_65#_M1019_g
+ N_A_149_65#_M1016_g N_A_149_65#_c_471_n N_A_149_65#_c_478_n
+ N_A_149_65#_c_472_n N_A_149_65#_c_473_n N_A_149_65#_c_506_n
+ N_A_149_65#_c_474_n N_A_149_65#_c_475_n PM_SKY130_FD_SC_LP__XOR2_2%A_149_65#
x_PM_SKY130_FD_SC_LP__XOR2_2%VPWR N_VPWR_M1001_s N_VPWR_M1015_s N_VPWR_M1006_d
+ N_VPWR_M1017_d N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n
+ N_VPWR_c_587_n VPWR N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n
+ N_VPWR_c_582_n N_VPWR_c_592_n N_VPWR_c_593_n N_VPWR_c_594_n
+ PM_SKY130_FD_SC_LP__XOR2_2%VPWR
x_PM_SKY130_FD_SC_LP__XOR2_2%A_149_367# N_A_149_367#_M1001_d
+ N_A_149_367#_M1014_d N_A_149_367#_c_684_n N_A_149_367#_c_671_n
+ N_A_149_367#_c_673_n N_A_149_367#_c_675_n
+ PM_SKY130_FD_SC_LP__XOR2_2%A_149_367#
x_PM_SKY130_FD_SC_LP__XOR2_2%A_532_367# N_A_532_367#_M1002_s
+ N_A_532_367#_M1016_s N_A_532_367#_M1005_s N_A_532_367#_M1013_s
+ N_A_532_367#_c_704_n N_A_532_367#_c_690_n N_A_532_367#_c_691_n
+ N_A_532_367#_c_698_n PM_SKY130_FD_SC_LP__XOR2_2%A_532_367#
x_PM_SKY130_FD_SC_LP__XOR2_2%X N_X_M1007_s N_X_M1012_s N_X_M1002_d N_X_c_779_n
+ N_X_c_741_n N_X_c_737_n N_X_c_786_n N_X_c_732_n N_X_c_753_n N_X_c_733_n X X X
+ X N_X_c_735_n X PM_SKY130_FD_SC_LP__XOR2_2%X
x_PM_SKY130_FD_SC_LP__XOR2_2%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_M1004_d
+ N_VGND_M1019_d N_VGND_M1010_s N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n
+ N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n
+ N_VGND_c_834_n N_VGND_c_835_n VGND N_VGND_c_836_n N_VGND_c_837_n
+ N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n PM_SKY130_FD_SC_LP__XOR2_2%VGND
x_PM_SKY130_FD_SC_LP__XOR2_2%A_814_65# N_A_814_65#_M1008_d N_A_814_65#_M1018_d
+ N_A_814_65#_c_899_n N_A_814_65#_c_900_n N_A_814_65#_c_901_n
+ N_A_814_65#_c_902_n PM_SKY130_FD_SC_LP__XOR2_2%A_814_65#
cc_1 VNB N_A_M1001_g 0.00374192f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.465
cc_2 VNB N_A_M1004_g 0.0248283f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=0.745
cc_3 VNB N_A_M1006_g 0.00224118f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=2.465
cc_4 VNB N_A_M1010_g 0.0257258f $X=-0.19 $Y=-0.245 $X2=5.675 $Y2=0.745
cc_5 VNB N_A_c_106_n 0.00727355f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.345
cc_6 VNB N_A_c_107_n 5.32246e-19 $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.95
cc_7 VNB N_A_c_108_n 0.0018089f $X=-0.19 $Y=-0.245 $X2=3.83 $Y2=1.355
cc_8 VNB N_A_c_109_n 2.10274e-19 $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.92
cc_9 VNB N_A_c_110_n 0.0362889f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.44
cc_10 VNB N_A_c_111_n 0.0133684f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.475
cc_11 VNB N_A_c_112_n 0.0303871f $X=-0.19 $Y=-0.245 $X2=3.905 $Y2=1.44
cc_12 VNB N_A_c_113_n 0.00383851f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.48
cc_13 VNB N_A_c_114_n 0.0188663f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.275
cc_14 VNB N_A_c_115_n 0.0019759f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=1.51
cc_15 VNB N_A_c_116_n 0.0314837f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.51
cc_16 VNB N_A_c_117_n 0.0186299f $X=-0.19 $Y=-0.245 $X2=3.905 $Y2=1.275
cc_17 VNB N_A_c_118_n 0.0320123f $X=-0.19 $Y=-0.245 $X2=5.675 $Y2=1.51
cc_18 VNB N_B_M1009_g 0.0224834f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.745
cc_19 VNB N_B_M1011_g 0.0248218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_M1012_g 0.0200844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_M1018_g 0.0227706f $X=-0.19 $Y=-0.245 $X2=5.675 $Y2=1.345
cc_22 VNB N_B_c_328_n 0.0118726f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=0.7
cc_23 VNB N_B_c_329_n 0.00353998f $X=-0.19 $Y=-0.245 $X2=5.56 $Y2=1.51
cc_24 VNB N_B_c_330_n 0.0387657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_c_331_n 0.0409613f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.035
cc_26 VNB N_A_149_65#_c_467_n 0.0185761f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.465
cc_27 VNB N_A_149_65#_M1002_g 0.00246517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_149_65#_c_469_n 0.0179134f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=2.465
cc_29 VNB N_A_149_65#_M1016_g 0.00210882f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=0.745
cc_30 VNB N_A_149_65#_c_471_n 0.0153512f $X=-0.19 $Y=-0.245 $X2=5.47 $Y2=2.465
cc_31 VNB N_A_149_65#_c_472_n 0.00320885f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=0.7
cc_32 VNB N_A_149_65#_c_473_n 5.9194e-19 $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.605
cc_33 VNB N_A_149_65#_c_474_n 0.00221753f $X=-0.19 $Y=-0.245 $X2=5.56 $Y2=1.51
cc_34 VNB N_A_149_65#_c_475_n 0.0588482f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.44
cc_35 VNB N_VPWR_c_582_n 0.263193f $X=-0.19 $Y=-0.245 $X2=5.56 $Y2=1.51
cc_36 VNB N_X_c_732_n 0.0114385f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=2.465
cc_37 VNB N_X_c_733_n 0.00137526f $X=-0.19 $Y=-0.245 $X2=5.47 $Y2=2.465
cc_38 VNB X 0.00515492f $X=-0.19 $Y=-0.245 $X2=5.675 $Y2=1.345
cc_39 VNB N_X_c_735_n 0.0094505f $X=-0.19 $Y=-0.245 $X2=3.83 $Y2=1.355
cc_40 VNB X 0.0215336f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.92
cc_41 VNB N_VGND_c_826_n 0.0147344f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=1.605
cc_42 VNB N_VGND_c_827_n 0.0157501f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=2.465
cc_43 VNB N_VGND_c_828_n 0.00736959f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=0.745
cc_44 VNB N_VGND_c_829_n 0.00738861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_830_n 0.0196648f $X=-0.19 $Y=-0.245 $X2=5.675 $Y2=0.745
cc_46 VNB N_VGND_c_831_n 0.00712408f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.345
cc_47 VNB N_VGND_c_832_n 0.0122131f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.7
cc_48 VNB N_VGND_c_833_n 0.0332136f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.95
cc_49 VNB N_VGND_c_834_n 0.0191207f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.605
cc_50 VNB N_VGND_c_835_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.92
cc_51 VNB N_VGND_c_836_n 0.0249686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_837_n 0.0462642f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.44
cc_53 VNB N_VGND_c_838_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.95
cc_54 VNB N_VGND_c_839_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_840_n 0.338819f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.51
cc_56 VNB N_A_814_65#_c_899_n 0.00372208f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.465
cc_57 VNB N_A_814_65#_c_900_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_814_65#_c_901_n 0.00221542f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.345
cc_59 VNB N_A_814_65#_c_902_n 0.00526341f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=0.745
cc_60 VPB N_A_M1001_g 0.0258373f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.465
cc_61 VPB N_A_M1015_g 0.0225964f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=2.465
cc_62 VPB N_A_M1006_g 0.0206556f $X=-0.19 $Y=1.655 $X2=3.86 $Y2=2.465
cc_63 VPB N_A_M1013_g 0.0250023f $X=-0.19 $Y=1.655 $X2=5.47 $Y2=2.465
cc_64 VPB N_A_c_107_n 0.00115549f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.95
cc_65 VPB N_A_c_109_n 0.00114164f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.92
cc_66 VPB N_A_c_125_n 0.00148678f $X=-0.19 $Y=1.655 $X2=5.56 $Y2=1.51
cc_67 VPB N_A_c_115_n 0.00102974f $X=-0.19 $Y=1.655 $X2=2.17 $Y2=1.51
cc_68 VPB N_A_c_116_n 0.0106399f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=1.51
cc_69 VPB N_A_c_118_n 0.00776019f $X=-0.19 $Y=1.655 $X2=5.675 $Y2=1.51
cc_70 VPB N_B_M1000_g 0.018015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_B_M1014_g 0.0188281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B_M1005_g 0.0197559f $X=-0.19 $Y=1.655 $X2=5.47 $Y2=1.675
cc_73 VPB N_B_M1017_g 0.0203206f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=0.785
cc_74 VPB N_B_c_328_n 0.0157315f $X=-0.19 $Y=1.655 $X2=3.74 $Y2=0.7
cc_75 VPB N_B_c_337_n 0.00122347f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.7
cc_76 VPB B 0.00170258f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.605
cc_77 VPB N_B_c_329_n 0.00266994f $X=-0.19 $Y=1.655 $X2=5.56 $Y2=1.51
cc_78 VPB N_B_c_330_n 0.00946488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_B_c_341_n 0.00273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_B_c_331_n 0.00766463f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.035
cc_81 VPB N_A_149_65#_M1002_g 0.0237231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_149_65#_M1016_g 0.0189711f $X=-0.19 $Y=1.655 $X2=3.995 $Y2=0.745
cc_83 VPB N_A_149_65#_c_478_n 0.0114428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_149_65#_c_473_n 0.00907442f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.605
cc_85 VPB N_VPWR_c_583_n 0.0234637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_584_n 0.0432749f $X=-0.19 $Y=1.655 $X2=3.86 $Y2=2.465
cc_87 VPB N_VPWR_c_585_n 0.00747655f $X=-0.19 $Y=1.655 $X2=3.995 $Y2=0.745
cc_88 VPB N_VPWR_c_586_n 0.0183997f $X=-0.19 $Y=1.655 $X2=5.47 $Y2=1.675
cc_89 VPB N_VPWR_c_587_n 0.00712965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_588_n 0.0339128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_589_n 0.0371113f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.605
cc_92 VPB N_VPWR_c_590_n 0.0281855f $X=-0.19 $Y=1.655 $X2=5.56 $Y2=1.51
cc_93 VPB N_VPWR_c_582_n 0.0717263f $X=-0.19 $Y=1.655 $X2=5.56 $Y2=1.51
cc_94 VPB N_VPWR_c_592_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.44
cc_95 VPB N_VPWR_c_593_n 0.0109593f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.035
cc_96 VPB N_VPWR_c_594_n 0.0109593f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.95
cc_97 VPB N_A_532_367#_c_690_n 0.00468671f $X=-0.19 $Y=1.655 $X2=2.35 $Y2=0.745
cc_98 VPB N_A_532_367#_c_691_n 0.00792372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_X_c_737_n 0.0243528f $X=-0.19 $Y=1.655 $X2=3.86 $Y2=1.605
cc_100 VPB N_X_c_733_n 0.00151682f $X=-0.19 $Y=1.655 $X2=5.47 $Y2=2.465
cc_101 VPB X 0.0324375f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.92
cc_102 N_A_c_106_n N_B_M1009_g 2.96382e-19 $X=0.455 $Y=1.345 $X2=0 $Y2=0
cc_103 N_A_c_130_p N_B_M1009_g 0.0124018f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_104 N_A_c_114_n N_B_M1009_g 0.02938f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_105 N_A_M1001_g N_B_M1000_g 0.02938f $X=0.67 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_c_107_n N_B_M1000_g 0.00345572f $X=0.76 $Y=1.95 $X2=0 $Y2=0
cc_107 A N_B_M1000_g 0.0149583f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_108 N_A_c_115_n N_B_M1000_g 8.97149e-19 $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A_M1015_g N_B_M1014_g 0.0428497f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_110 A N_B_M1014_g 0.00833389f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_111 N_A_c_115_n N_B_M1014_g 0.0106233f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_112 N_A_M1004_g N_B_M1011_g 0.0293466f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_113 N_A_c_130_p N_B_M1011_g 0.0134264f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_114 N_A_c_108_n N_B_M1012_g 3.2667e-19 $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_115 N_A_c_117_n N_B_M1012_g 0.0199484f $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_116 N_A_M1006_g N_B_M1005_g 0.0407879f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_c_109_n N_B_M1005_g 0.00338052f $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_118 N_A_c_145_p N_B_M1005_g 0.0111311f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_119 N_A_M1010_g N_B_M1018_g 0.00891267f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_120 N_A_M1013_g N_B_M1017_g 0.026067f $X=5.47 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_c_145_p N_B_M1017_g 0.0111875f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_122 N_A_M1006_g N_B_c_328_n 0.00242047f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_c_108_n N_B_c_328_n 7.00442e-19 $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_124 N_A_c_109_n N_B_c_328_n 0.0097379f $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_125 N_A_c_145_p N_B_c_328_n 0.0105813f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_126 N_A_c_112_n N_B_c_328_n 5.56753e-19 $X=3.905 $Y=1.44 $X2=0 $Y2=0
cc_127 N_A_c_113_n N_B_c_328_n 0.0121277f $X=3.985 $Y=1.48 $X2=0 $Y2=0
cc_128 A N_B_c_328_n 0.00691405f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_129 N_A_c_115_n N_B_c_328_n 0.0398386f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A_c_116_n N_B_c_328_n 0.00264334f $X=2.35 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A_c_107_n N_B_c_337_n 0.00115434f $X=0.76 $Y=1.95 $X2=0 $Y2=0
cc_132 N_A_c_111_n N_B_c_337_n 3.96424e-19 $X=0.76 $Y=1.475 $X2=0 $Y2=0
cc_133 A N_B_c_337_n 0.00216454f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_134 N_A_c_115_n N_B_c_337_n 5.78644e-19 $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A_c_109_n B 0.00120221f $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_136 N_A_c_145_p B 0.00776137f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_137 N_A_c_113_n B 2.41172e-19 $X=3.985 $Y=1.48 $X2=0 $Y2=0
cc_138 N_A_M1001_g N_B_c_329_n 5.04626e-19 $X=0.67 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_c_107_n N_B_c_329_n 0.0129695f $X=0.76 $Y=1.95 $X2=0 $Y2=0
cc_140 N_A_c_110_n N_B_c_329_n 7.38433e-19 $X=0.58 $Y=1.44 $X2=0 $Y2=0
cc_141 N_A_c_111_n N_B_c_329_n 0.0221328f $X=0.76 $Y=1.475 $X2=0 $Y2=0
cc_142 A N_B_c_329_n 0.0244787f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_143 N_A_c_115_n N_B_c_329_n 0.0328897f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A_c_107_n N_B_c_330_n 5.37505e-19 $X=0.76 $Y=1.95 $X2=0 $Y2=0
cc_145 N_A_c_110_n N_B_c_330_n 0.02938f $X=0.58 $Y=1.44 $X2=0 $Y2=0
cc_146 N_A_c_111_n N_B_c_330_n 9.35219e-19 $X=0.76 $Y=1.475 $X2=0 $Y2=0
cc_147 A N_B_c_330_n 5.38132e-19 $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_148 N_A_c_115_n N_B_c_330_n 0.0184647f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A_c_116_n N_B_c_330_n 0.0215485f $X=2.35 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A_M1006_g N_B_c_341_n 3.0878e-19 $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_c_109_n N_B_c_341_n 0.00814297f $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_152 N_A_c_145_p N_B_c_341_n 0.0405277f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_153 N_A_c_125_n N_B_c_341_n 0.0122729f $X=5.56 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A_c_112_n N_B_c_341_n 2.44541e-19 $X=3.905 $Y=1.44 $X2=0 $Y2=0
cc_155 N_A_c_113_n N_B_c_341_n 0.0120802f $X=3.985 $Y=1.48 $X2=0 $Y2=0
cc_156 N_A_c_118_n N_B_c_341_n 0.00138908f $X=5.675 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A_M1006_g N_B_c_331_n 0.00259342f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_c_109_n N_B_c_331_n 3.75466e-19 $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_159 N_A_c_145_p N_B_c_331_n 9.81766e-19 $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_160 N_A_c_125_n N_B_c_331_n 0.0024897f $X=5.56 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A_c_112_n N_B_c_331_n 0.0168662f $X=3.905 $Y=1.44 $X2=0 $Y2=0
cc_162 N_A_c_113_n N_B_c_331_n 0.00120799f $X=3.985 $Y=1.48 $X2=0 $Y2=0
cc_163 N_A_c_118_n N_B_c_331_n 0.026067f $X=5.675 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A_c_130_p N_A_149_65#_M1003_s 0.00459188f $X=3.74 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_c_130_p N_A_149_65#_M1011_s 0.0121022f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_166 A N_A_149_65#_M1000_s 0.00319681f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_167 N_A_M1004_g N_A_149_65#_c_467_n 0.0245142f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_168 N_A_c_130_p N_A_149_65#_c_467_n 0.0140376f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_169 N_A_c_116_n N_A_149_65#_M1002_g 0.00177691f $X=2.35 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A_c_130_p N_A_149_65#_c_469_n 0.0154158f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_171 N_A_c_108_n N_A_149_65#_c_469_n 0.00593847f $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_172 N_A_c_117_n N_A_149_65#_c_469_n 0.0230469f $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_173 N_A_M1006_g N_A_149_65#_M1016_g 0.0561421f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_c_109_n N_A_149_65#_M1016_g 9.7149e-19 $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_175 N_A_c_202_p N_A_149_65#_M1016_g 5.0656e-19 $X=4.07 $Y=2.005 $X2=0 $Y2=0
cc_176 N_A_M1004_g N_A_149_65#_c_471_n 0.0146326f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_177 N_A_c_106_n N_A_149_65#_c_471_n 0.00905947f $X=0.455 $Y=1.345 $X2=0 $Y2=0
cc_178 N_A_c_130_p N_A_149_65#_c_471_n 0.115256f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_179 N_A_c_111_n N_A_149_65#_c_471_n 0.00971729f $X=0.76 $Y=1.475 $X2=0 $Y2=0
cc_180 N_A_c_114_n N_A_149_65#_c_471_n 0.00316042f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_181 N_A_c_115_n N_A_149_65#_c_471_n 0.0574882f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_c_116_n N_A_149_65#_c_471_n 0.00735745f $X=2.35 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A_M1015_g N_A_149_65#_c_478_n 0.016636f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_184 A N_A_149_65#_c_478_n 0.0532369f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_185 N_A_c_116_n N_A_149_65#_c_478_n 0.00219802f $X=2.35 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A_M1004_g N_A_149_65#_c_472_n 0.00366784f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A_M1015_g N_A_149_65#_c_473_n 0.00645439f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_c_115_n N_A_149_65#_c_473_n 0.0368633f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_189 N_A_c_116_n N_A_149_65#_c_473_n 5.7708e-19 $X=2.35 $Y=1.51 $X2=0 $Y2=0
cc_190 A N_A_149_65#_c_506_n 0.0123465f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_191 N_A_M1004_g N_A_149_65#_c_474_n 0.00256611f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_192 N_A_c_130_p N_A_149_65#_c_474_n 0.00840781f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_193 N_A_c_115_n N_A_149_65#_c_474_n 0.0200717f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A_M1004_g N_A_149_65#_c_475_n 0.0145726f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_195 N_A_c_130_p N_A_149_65#_c_475_n 0.0033865f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_196 N_A_c_108_n N_A_149_65#_c_475_n 3.63824e-19 $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_197 N_A_c_112_n N_A_149_65#_c_475_n 0.0191885f $X=3.905 $Y=1.44 $X2=0 $Y2=0
cc_198 N_A_c_113_n N_A_149_65#_c_475_n 0.00112447f $X=3.985 $Y=1.48 $X2=0 $Y2=0
cc_199 N_A_c_115_n N_A_149_65#_c_475_n 2.19001e-19 $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A_c_115_n N_VPWR_M1015_s 0.00517725f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A_c_109_n N_VPWR_M1006_d 0.00108503f $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_202 N_A_c_145_p N_VPWR_M1006_d 0.00645472f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_203 N_A_c_202_p N_VPWR_M1006_d 8.45435e-19 $X=4.07 $Y=2.005 $X2=0 $Y2=0
cc_204 N_A_c_145_p N_VPWR_M1017_d 0.0111229f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_205 N_A_M1001_g N_VPWR_c_583_n 0.00608886f $X=0.67 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_c_107_n N_VPWR_c_583_n 0.00939472f $X=0.76 $Y=1.95 $X2=0 $Y2=0
cc_207 N_A_c_110_n N_VPWR_c_583_n 0.00202522f $X=0.58 $Y=1.44 $X2=0 $Y2=0
cc_208 N_A_c_111_n N_VPWR_c_583_n 0.00951325f $X=0.76 $Y=1.475 $X2=0 $Y2=0
cc_209 N_A_c_236_p N_VPWR_c_583_n 0.0137304f $X=0.845 $Y=2.035 $X2=0 $Y2=0
cc_210 N_A_M1001_g N_VPWR_c_584_n 0.014552f $X=0.67 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_M1015_g N_VPWR_c_585_n 0.0140988f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_M1001_g N_VPWR_c_587_n 0.00303312f $X=0.67 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_c_110_n N_VPWR_c_587_n 0.00154266f $X=0.58 $Y=1.44 $X2=0 $Y2=0
cc_214 N_A_M1001_g N_VPWR_c_588_n 0.00486043f $X=0.67 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_M1015_g N_VPWR_c_588_n 0.00486043f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_M1006_g N_VPWR_c_589_n 0.00404333f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_M1013_g N_VPWR_c_590_n 0.00413624f $X=5.47 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_M1001_g N_VPWR_c_582_n 0.0082726f $X=0.67 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A_M1015_g N_VPWR_c_582_n 0.00859951f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A_M1006_g N_VPWR_c_582_n 0.00607537f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A_M1013_g N_VPWR_c_582_n 0.00732249f $X=5.47 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A_M1006_g N_VPWR_c_593_n 0.00408156f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A_M1013_g N_VPWR_c_594_n 0.00408156f $X=5.47 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_c_107_n N_A_149_367#_M1001_d 0.00133118f $X=0.76 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A_c_236_p N_A_149_367#_M1001_d 4.60859e-19 $X=0.845 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_226 A N_A_149_367#_M1001_d 0.00595186f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_227 N_A_c_115_n N_A_149_367#_M1014_d 0.00299302f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_c_236_p N_A_149_367#_c_671_n 0.00375541f $X=0.845 $Y=2.035 $X2=0
+ $Y2=0
cc_229 A N_A_149_367#_c_671_n 0.00997062f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_230 N_A_c_145_p N_A_532_367#_M1005_s 0.00321722f $X=5.395 $Y=2.005 $X2=0
+ $Y2=0
cc_231 N_A_c_145_p N_A_532_367#_M1013_s 0.00323899f $X=5.395 $Y=2.005 $X2=0
+ $Y2=0
cc_232 N_A_c_125_n N_A_532_367#_M1013_s 9.1358e-19 $X=5.56 $Y=1.51 $X2=0 $Y2=0
cc_233 N_A_M1015_g N_A_532_367#_c_690_n 0.00111902f $X=2.05 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A_M1006_g N_A_532_367#_c_691_n 0.0089268f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A_M1013_g N_A_532_367#_c_691_n 0.0101574f $X=5.47 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_M1006_g N_A_532_367#_c_698_n 0.00727308f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_c_130_p N_X_M1007_s 0.00447029f $X=3.74 $Y=0.7 $X2=-0.19 $Y2=-0.245
cc_238 N_A_c_202_p N_X_c_741_n 0.00540651f $X=4.07 $Y=2.005 $X2=0 $Y2=0
cc_239 N_A_M1006_g N_X_c_737_n 0.0127656f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_M1013_g N_X_c_737_n 0.0131006f $X=5.47 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A_c_145_p N_X_c_737_n 0.0939851f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_242 N_A_c_202_p N_X_c_737_n 0.00842766f $X=4.07 $Y=2.005 $X2=0 $Y2=0
cc_243 N_A_c_112_n N_X_c_737_n 3.02919e-19 $X=3.905 $Y=1.44 $X2=0 $Y2=0
cc_244 N_A_c_113_n N_X_c_737_n 0.00136355f $X=3.985 $Y=1.48 $X2=0 $Y2=0
cc_245 N_A_c_118_n N_X_c_737_n 0.00116495f $X=5.675 $Y=1.51 $X2=0 $Y2=0
cc_246 N_A_M1010_g N_X_c_732_n 0.0179813f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_247 N_A_c_145_p N_X_c_732_n 0.0066003f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_248 N_A_c_125_n N_X_c_732_n 0.0257317f $X=5.56 $Y=1.51 $X2=0 $Y2=0
cc_249 N_A_c_118_n N_X_c_732_n 0.00564371f $X=5.675 $Y=1.51 $X2=0 $Y2=0
cc_250 N_A_c_130_p N_X_c_753_n 0.0173168f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_251 N_A_c_108_n N_X_c_753_n 0.0085209f $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_252 N_A_M1006_g N_X_c_733_n 0.00227286f $X=3.86 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A_c_108_n N_X_c_733_n 0.00768519f $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_254 N_A_c_109_n N_X_c_733_n 0.00698706f $X=3.985 $Y=1.92 $X2=0 $Y2=0
cc_255 N_A_c_112_n N_X_c_733_n 5.20499e-19 $X=3.905 $Y=1.44 $X2=0 $Y2=0
cc_256 N_A_c_113_n N_X_c_733_n 0.00960929f $X=3.985 $Y=1.48 $X2=0 $Y2=0
cc_257 N_A_M1010_g X 0.0031541f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_258 N_A_c_108_n X 0.00194307f $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_259 N_A_c_145_p X 0.00428642f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_260 N_A_c_117_n X 3.42363e-19 $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_261 N_A_M1013_g X 0.00704416f $X=5.47 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A_M1010_g X 0.0126736f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_263 N_A_c_145_p X 0.0144849f $X=5.395 $Y=2.005 $X2=0 $Y2=0
cc_264 N_A_c_125_n X 0.0400605f $X=5.56 $Y=1.51 $X2=0 $Y2=0
cc_265 N_A_c_106_n N_VGND_M1003_d 0.0161054f $X=0.455 $Y=1.345 $X2=-0.19
+ $Y2=-0.245
cc_266 N_A_c_293_p N_VGND_M1003_d 0.00995521f $X=0.54 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_267 N_A_c_130_p N_VGND_M1009_d 0.0072714f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_268 N_A_c_130_p N_VGND_M1004_d 0.00953252f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_269 N_A_c_130_p N_VGND_M1019_d 0.012958f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_270 N_A_c_108_n N_VGND_M1019_d 0.00667733f $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_271 N_A_c_293_p N_VGND_c_827_n 0.0128817f $X=0.54 $Y=0.7 $X2=0 $Y2=0
cc_272 N_A_c_114_n N_VGND_c_827_n 0.00995887f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_273 N_A_c_130_p N_VGND_c_828_n 0.0246925f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_274 N_A_M1004_g N_VGND_c_829_n 0.0043151f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_275 N_A_c_130_p N_VGND_c_829_n 0.0247682f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_276 N_A_c_130_p N_VGND_c_830_n 0.0110801f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_277 N_A_c_130_p N_VGND_c_831_n 0.0256321f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_278 N_A_c_117_n N_VGND_c_831_n 0.00292562f $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_279 N_A_M1010_g N_VGND_c_833_n 0.0150025f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_280 N_A_c_130_p N_VGND_c_834_n 0.0104671f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_281 N_A_c_293_p N_VGND_c_834_n 2.72161e-19 $X=0.54 $Y=0.7 $X2=0 $Y2=0
cc_282 N_A_c_114_n N_VGND_c_834_n 0.00353682f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_283 N_A_M1004_g N_VGND_c_836_n 0.00353682f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_284 N_A_c_130_p N_VGND_c_836_n 0.0146574f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_285 N_A_M1010_g N_VGND_c_837_n 0.00466675f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_286 N_A_c_117_n N_VGND_c_837_n 0.00499542f $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_287 N_A_M1004_g N_VGND_c_840_n 0.00515141f $X=2.35 $Y=0.745 $X2=0 $Y2=0
cc_288 N_A_M1010_g N_VGND_c_840_n 0.00950445f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_289 N_A_c_130_p N_VGND_c_840_n 0.0698553f $X=3.74 $Y=0.7 $X2=0 $Y2=0
cc_290 N_A_c_293_p N_VGND_c_840_n 0.00130788f $X=0.54 $Y=0.7 $X2=0 $Y2=0
cc_291 N_A_c_114_n N_VGND_c_840_n 0.00525866f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_292 N_A_c_117_n N_VGND_c_840_n 0.00995623f $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_293 N_A_c_108_n N_A_814_65#_c_899_n 0.00146187f $X=3.83 $Y=1.355 $X2=0 $Y2=0
cc_294 N_A_c_117_n N_A_814_65#_c_899_n 9.65679e-19 $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_295 N_A_c_117_n N_A_814_65#_c_901_n 6.87828e-19 $X=3.905 $Y=1.275 $X2=0 $Y2=0
cc_296 N_A_M1010_g N_A_814_65#_c_902_n 0.00884027f $X=5.675 $Y=0.745 $X2=0 $Y2=0
cc_297 N_B_c_328_n N_A_149_65#_M1002_g 0.00801352f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_298 N_B_c_328_n N_A_149_65#_M1016_g 0.00267139f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_299 N_B_M1009_g N_A_149_65#_c_471_n 0.010908f $X=1.1 $Y=0.745 $X2=0 $Y2=0
cc_300 N_B_M1011_g N_A_149_65#_c_471_n 0.0147286f $X=1.69 $Y=0.745 $X2=0 $Y2=0
cc_301 N_B_c_328_n N_A_149_65#_c_471_n 0.0157971f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_302 N_B_c_337_n N_A_149_65#_c_471_n 0.00136003f $X=1.345 $Y=1.665 $X2=0 $Y2=0
cc_303 N_B_c_329_n N_A_149_65#_c_471_n 0.0300884f $X=1.33 $Y=1.51 $X2=0 $Y2=0
cc_304 N_B_c_330_n N_A_149_65#_c_471_n 0.00543592f $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_305 N_B_M1014_g N_A_149_65#_c_478_n 0.00970081f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_306 N_B_c_328_n N_A_149_65#_c_478_n 0.00873558f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_307 N_B_c_330_n N_A_149_65#_c_478_n 3.96656e-19 $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_308 N_B_c_328_n N_A_149_65#_c_472_n 6.17318e-19 $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_309 N_B_c_328_n N_A_149_65#_c_473_n 0.0157868f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_310 N_B_c_328_n N_A_149_65#_c_474_n 0.0231867f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_311 N_B_c_328_n N_A_149_65#_c_475_n 0.0100322f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_312 N_B_M1000_g N_VPWR_c_584_n 0.00110057f $X=1.1 $Y=2.465 $X2=0 $Y2=0
cc_313 N_B_M1014_g N_VPWR_c_585_n 0.00116113f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_314 N_B_M1005_g N_VPWR_c_586_n 0.00413624f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_315 N_B_M1017_g N_VPWR_c_586_n 0.00413624f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_316 N_B_M1000_g N_VPWR_c_588_n 0.00357877f $X=1.1 $Y=2.465 $X2=0 $Y2=0
cc_317 N_B_M1014_g N_VPWR_c_588_n 0.00359389f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_318 N_B_M1000_g N_VPWR_c_582_n 0.00537654f $X=1.1 $Y=2.465 $X2=0 $Y2=0
cc_319 N_B_M1014_g N_VPWR_c_582_n 0.00562094f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_320 N_B_M1005_g N_VPWR_c_582_n 0.00611928f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_321 N_B_M1017_g N_VPWR_c_582_n 0.00611928f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_322 N_B_M1005_g N_VPWR_c_593_n 0.00408156f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_323 N_B_M1017_g N_VPWR_c_594_n 0.00408156f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_324 N_B_M1000_g N_A_149_367#_c_673_n 0.0153414f $X=1.1 $Y=2.465 $X2=0 $Y2=0
cc_325 N_B_M1014_g N_A_149_367#_c_673_n 0.0119405f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_326 N_B_M1000_g N_A_149_367#_c_675_n 5.51056e-19 $X=1.1 $Y=2.465 $X2=0 $Y2=0
cc_327 N_B_M1014_g N_A_149_367#_c_675_n 0.00537498f $X=1.53 $Y=2.465 $X2=0 $Y2=0
cc_328 N_B_M1005_g N_A_532_367#_c_691_n 0.0101916f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_329 N_B_M1017_g N_A_532_367#_c_691_n 0.0101574f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_330 N_B_M1005_g N_A_532_367#_c_698_n 7.88281e-19 $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_331 N_B_c_328_n N_X_c_741_n 0.00856393f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_332 N_B_M1005_g N_X_c_737_n 0.0112087f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_333 N_B_M1017_g N_X_c_737_n 0.0111936f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_334 N_B_c_328_n N_X_c_737_n 0.0146506f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_335 N_B_c_328_n N_X_c_753_n 0.00619887f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_336 N_B_c_328_n N_X_c_733_n 0.0202214f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_337 N_B_M1012_g X 0.00877957f $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_338 N_B_M1018_g X 0.0196063f $X=4.88 $Y=0.745 $X2=0 $Y2=0
cc_339 B X 0.00139926f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_340 N_B_c_341_n X 0.0379323f $X=4.79 $Y=1.51 $X2=0 $Y2=0
cc_341 N_B_c_331_n X 0.00326418f $X=4.88 $Y=1.51 $X2=0 $Y2=0
cc_342 N_B_M1009_g N_VGND_c_828_n 0.00421885f $X=1.1 $Y=0.745 $X2=0 $Y2=0
cc_343 N_B_M1011_g N_VGND_c_828_n 0.00421885f $X=1.69 $Y=0.745 $X2=0 $Y2=0
cc_344 N_B_M1009_g N_VGND_c_834_n 0.00353682f $X=1.1 $Y=0.745 $X2=0 $Y2=0
cc_345 N_B_M1011_g N_VGND_c_836_n 0.00353682f $X=1.69 $Y=0.745 $X2=0 $Y2=0
cc_346 N_B_M1012_g N_VGND_c_837_n 0.00302501f $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_347 N_B_M1018_g N_VGND_c_837_n 0.00302501f $X=4.88 $Y=0.745 $X2=0 $Y2=0
cc_348 N_B_M1009_g N_VGND_c_840_n 0.00495111f $X=1.1 $Y=0.745 $X2=0 $Y2=0
cc_349 N_B_M1011_g N_VGND_c_840_n 0.0051267f $X=1.69 $Y=0.745 $X2=0 $Y2=0
cc_350 N_B_M1012_g N_VGND_c_840_n 0.00438099f $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_351 N_B_M1018_g N_VGND_c_840_n 0.00463014f $X=4.88 $Y=0.745 $X2=0 $Y2=0
cc_352 N_B_M1012_g N_A_814_65#_c_899_n 9.16006e-19 $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_353 N_B_c_328_n N_A_814_65#_c_899_n 0.00822718f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_354 N_B_c_341_n N_A_814_65#_c_899_n 0.00109722f $X=4.79 $Y=1.51 $X2=0 $Y2=0
cc_355 N_B_c_331_n N_A_814_65#_c_899_n 4.86925e-19 $X=4.88 $Y=1.51 $X2=0 $Y2=0
cc_356 N_B_M1012_g N_A_814_65#_c_900_n 0.0119553f $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_357 N_B_M1018_g N_A_814_65#_c_900_n 0.00996097f $X=4.88 $Y=0.745 $X2=0 $Y2=0
cc_358 N_B_M1018_g N_A_814_65#_c_902_n 0.00178673f $X=4.88 $Y=0.745 $X2=0 $Y2=0
cc_359 N_A_149_65#_c_478_n N_VPWR_M1015_s 0.00494748f $X=2.53 $Y=2.375 $X2=0
+ $Y2=0
cc_360 N_A_149_65#_M1002_g N_VPWR_c_585_n 0.00338413f $X=3 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A_149_65#_c_478_n N_VPWR_c_585_n 0.0220026f $X=2.53 $Y=2.375 $X2=0
+ $Y2=0
cc_362 N_A_149_65#_M1002_g N_VPWR_c_589_n 0.00357668f $X=3 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A_149_65#_M1016_g N_VPWR_c_589_n 0.00357877f $X=3.43 $Y=2.465 $X2=0
+ $Y2=0
cc_364 N_A_149_65#_M1000_s N_VPWR_c_582_n 0.00225186f $X=1.175 $Y=1.835 $X2=0
+ $Y2=0
cc_365 N_A_149_65#_M1002_g N_VPWR_c_582_n 0.00682149f $X=3 $Y=2.465 $X2=0 $Y2=0
cc_366 N_A_149_65#_M1016_g N_VPWR_c_582_n 0.00544922f $X=3.43 $Y=2.465 $X2=0
+ $Y2=0
cc_367 N_A_149_65#_c_478_n N_A_149_367#_M1014_d 0.00540754f $X=2.53 $Y=2.375
+ $X2=0 $Y2=0
cc_368 N_A_149_65#_M1000_s N_A_149_367#_c_673_n 0.00337304f $X=1.175 $Y=1.835
+ $X2=0 $Y2=0
cc_369 N_A_149_65#_c_478_n N_A_149_367#_c_673_n 0.00583566f $X=2.53 $Y=2.375
+ $X2=0 $Y2=0
cc_370 N_A_149_65#_c_506_n N_A_149_367#_c_673_n 0.0126773f $X=1.31 $Y=2.375
+ $X2=0 $Y2=0
cc_371 N_A_149_65#_c_478_n N_A_149_367#_c_675_n 0.0203821f $X=2.53 $Y=2.375
+ $X2=0 $Y2=0
cc_372 N_A_149_65#_c_478_n N_A_532_367#_M1002_s 0.00291806f $X=2.53 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_373 N_A_149_65#_c_473_n N_A_532_367#_M1002_s 0.0062189f $X=2.615 $Y=2.29
+ $X2=-0.19 $Y2=-0.245
cc_374 N_A_149_65#_M1016_g N_A_532_367#_c_704_n 0.0168006f $X=3.43 $Y=2.465
+ $X2=0 $Y2=0
cc_375 N_A_149_65#_M1002_g N_A_532_367#_c_690_n 0.0230646f $X=3 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_A_149_65#_c_478_n N_A_532_367#_c_690_n 0.00708364f $X=2.53 $Y=2.375
+ $X2=0 $Y2=0
cc_377 N_A_149_65#_M1002_g N_X_c_779_n 0.00386807f $X=3 $Y=2.465 $X2=0 $Y2=0
cc_378 N_A_149_65#_M1016_g N_X_c_779_n 0.00453777f $X=3.43 $Y=2.465 $X2=0 $Y2=0
cc_379 N_A_149_65#_M1002_g N_X_c_741_n 0.00291561f $X=3 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A_149_65#_M1016_g N_X_c_741_n 0.00285008f $X=3.43 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A_149_65#_c_473_n N_X_c_741_n 0.0177543f $X=2.615 $Y=2.29 $X2=0 $Y2=0
cc_382 N_A_149_65#_c_475_n N_X_c_741_n 0.00156612f $X=3.43 $Y=1.44 $X2=0 $Y2=0
cc_383 N_A_149_65#_M1016_g N_X_c_737_n 0.00842512f $X=3.43 $Y=2.465 $X2=0 $Y2=0
cc_384 N_A_149_65#_M1002_g N_X_c_786_n 0.00293349f $X=3 $Y=2.465 $X2=0 $Y2=0
cc_385 N_A_149_65#_M1016_g N_X_c_786_n 7.17598e-19 $X=3.43 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A_149_65#_c_478_n N_X_c_786_n 0.00699722f $X=2.53 $Y=2.375 $X2=0 $Y2=0
cc_387 N_A_149_65#_c_473_n N_X_c_786_n 0.0013268f $X=2.615 $Y=2.29 $X2=0 $Y2=0
cc_388 N_A_149_65#_c_467_n N_X_c_753_n 0.0036641f $X=2.975 $Y=1.275 $X2=0 $Y2=0
cc_389 N_A_149_65#_c_469_n N_X_c_753_n 0.00417817f $X=3.405 $Y=1.275 $X2=0 $Y2=0
cc_390 N_A_149_65#_c_471_n N_X_c_753_n 0.0102683f $X=2.53 $Y=1.065 $X2=0 $Y2=0
cc_391 N_A_149_65#_c_474_n N_X_c_753_n 3.4131e-19 $X=2.865 $Y=1.44 $X2=0 $Y2=0
cc_392 N_A_149_65#_c_475_n N_X_c_753_n 0.00316943f $X=3.43 $Y=1.44 $X2=0 $Y2=0
cc_393 N_A_149_65#_c_467_n N_X_c_733_n 0.0010446f $X=2.975 $Y=1.275 $X2=0 $Y2=0
cc_394 N_A_149_65#_M1002_g N_X_c_733_n 0.00201605f $X=3 $Y=2.465 $X2=0 $Y2=0
cc_395 N_A_149_65#_c_469_n N_X_c_733_n 0.00275392f $X=3.405 $Y=1.275 $X2=0 $Y2=0
cc_396 N_A_149_65#_M1016_g N_X_c_733_n 0.00513291f $X=3.43 $Y=2.465 $X2=0 $Y2=0
cc_397 N_A_149_65#_c_471_n N_X_c_733_n 5.69824e-19 $X=2.53 $Y=1.065 $X2=0 $Y2=0
cc_398 N_A_149_65#_c_472_n N_X_c_733_n 0.00519301f $X=2.615 $Y=1.33 $X2=0 $Y2=0
cc_399 N_A_149_65#_c_473_n N_X_c_733_n 0.00646626f $X=2.615 $Y=2.29 $X2=0 $Y2=0
cc_400 N_A_149_65#_c_474_n N_X_c_733_n 0.0192725f $X=2.865 $Y=1.44 $X2=0 $Y2=0
cc_401 N_A_149_65#_c_475_n N_X_c_733_n 0.0159777f $X=3.43 $Y=1.44 $X2=0 $Y2=0
cc_402 N_A_149_65#_c_471_n N_VGND_M1009_d 0.00442708f $X=2.53 $Y=1.065 $X2=0
+ $Y2=0
cc_403 N_A_149_65#_c_471_n N_VGND_M1004_d 0.00577218f $X=2.53 $Y=1.065 $X2=0
+ $Y2=0
cc_404 N_A_149_65#_c_467_n N_VGND_c_829_n 0.00674628f $X=2.975 $Y=1.275 $X2=0
+ $Y2=0
cc_405 N_A_149_65#_c_467_n N_VGND_c_830_n 0.00353682f $X=2.975 $Y=1.275 $X2=0
+ $Y2=0
cc_406 N_A_149_65#_c_469_n N_VGND_c_830_n 0.00353682f $X=3.405 $Y=1.275 $X2=0
+ $Y2=0
cc_407 N_A_149_65#_c_469_n N_VGND_c_831_n 0.00421885f $X=3.405 $Y=1.275 $X2=0
+ $Y2=0
cc_408 N_A_149_65#_c_467_n N_VGND_c_840_n 0.00504448f $X=2.975 $Y=1.275 $X2=0
+ $Y2=0
cc_409 N_A_149_65#_c_469_n N_VGND_c_840_n 0.00494239f $X=3.405 $Y=1.275 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_582_n N_A_149_367#_M1001_d 0.00373407f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_411 N_VPWR_c_582_n N_A_149_367#_M1014_d 0.00457565f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_412 N_VPWR_c_588_n N_A_149_367#_c_684_n 0.0139427f $X=2.1 $Y=3.33 $X2=0 $Y2=0
cc_413 N_VPWR_c_582_n N_A_149_367#_c_684_n 0.00894187f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_414 N_VPWR_c_588_n N_A_149_367#_c_673_n 0.0337777f $X=2.1 $Y=3.33 $X2=0 $Y2=0
cc_415 N_VPWR_c_582_n N_A_149_367#_c_673_n 0.0206164f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_416 N_VPWR_c_588_n N_A_149_367#_c_675_n 0.0201338f $X=2.1 $Y=3.33 $X2=0 $Y2=0
cc_417 N_VPWR_c_582_n N_A_149_367#_c_675_n 0.0125965f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_c_582_n N_A_532_367#_M1002_s 0.00215962f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_419 N_VPWR_c_582_n N_A_532_367#_M1016_s 0.00225186f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_582_n N_A_532_367#_M1005_s 0.00296296f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_421 N_VPWR_c_582_n N_A_532_367#_M1013_s 0.00283281f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_422 N_VPWR_c_589_n N_A_532_367#_c_704_n 0.0353423f $X=3.99 $Y=3.33 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_582_n N_A_532_367#_c_704_n 0.0225965f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_424 N_VPWR_c_585_n N_A_532_367#_c_690_n 0.0363853f $X=2.265 $Y=2.755 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_589_n N_A_532_367#_c_690_n 0.0357549f $X=3.99 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_582_n N_A_532_367#_c_690_n 0.0217125f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_427 N_VPWR_M1006_d N_A_532_367#_c_691_n 0.00748372f $X=3.935 $Y=1.835 $X2=0
+ $Y2=0
cc_428 N_VPWR_M1017_d N_A_532_367#_c_691_n 0.00749438f $X=4.955 $Y=1.835 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_586_n N_A_532_367#_c_691_n 0.0119829f $X=5.01 $Y=3.33 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_589_n N_A_532_367#_c_691_n 0.00309909f $X=3.99 $Y=3.33 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_590_n N_A_532_367#_c_691_n 0.0094477f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_432 N_VPWR_c_582_n N_A_532_367#_c_691_n 0.0422512f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_433 N_VPWR_c_593_n N_A_532_367#_c_691_n 0.0242216f $X=4.155 $Y=3.025 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_594_n N_A_532_367#_c_691_n 0.0242216f $X=5.175 $Y=3.025 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_582_n N_X_M1002_d 0.00225177f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_436 N_VPWR_M1006_d N_X_c_737_n 0.00752182f $X=3.935 $Y=1.835 $X2=0 $Y2=0
cc_437 N_VPWR_M1017_d N_X_c_737_n 0.00769169f $X=4.955 $Y=1.835 $X2=0 $Y2=0
cc_438 N_A_532_367#_c_704_n N_X_M1002_d 0.00196301f $X=3.573 $Y=2.837 $X2=0
+ $Y2=0
cc_439 N_A_532_367#_c_690_n N_X_M1002_d 0.00144321f $X=3.202 $Y=2.837 $X2=0
+ $Y2=0
cc_440 N_A_532_367#_M1016_s N_X_c_737_n 0.00490421f $X=3.505 $Y=1.835 $X2=0
+ $Y2=0
cc_441 N_A_532_367#_M1005_s N_X_c_737_n 0.00341221f $X=4.525 $Y=1.835 $X2=0
+ $Y2=0
cc_442 N_A_532_367#_M1013_s N_X_c_737_n 0.00689165f $X=5.545 $Y=1.835 $X2=0
+ $Y2=0
cc_443 N_A_532_367#_c_704_n N_X_c_737_n 0.140173f $X=3.573 $Y=2.837 $X2=0 $Y2=0
cc_444 N_A_532_367#_c_704_n N_X_c_786_n 0.0103068f $X=3.573 $Y=2.837 $X2=0 $Y2=0
cc_445 N_A_532_367#_c_690_n N_X_c_786_n 0.00807896f $X=3.202 $Y=2.837 $X2=0
+ $Y2=0
cc_446 N_X_c_732_n N_VGND_M1010_s 9.24827e-19 $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_447 N_X_c_735_n N_VGND_M1010_s 0.00287472f $X=6.025 $Y=1.245 $X2=0 $Y2=0
cc_448 N_X_c_732_n N_VGND_c_833_n 0.00712308f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_449 N_X_c_735_n N_VGND_c_833_n 0.0207849f $X=6.025 $Y=1.245 $X2=0 $Y2=0
cc_450 N_X_c_732_n N_A_814_65#_M1018_d 0.00687105f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_451 X N_A_814_65#_M1018_d 0.00514876f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_452 X N_A_814_65#_c_899_n 0.0245772f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_453 N_X_M1012_s N_A_814_65#_c_900_n 0.00203037f $X=4.5 $Y=0.325 $X2=0 $Y2=0
cc_454 X N_A_814_65#_c_900_n 0.0210387f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_455 N_X_c_732_n N_A_814_65#_c_902_n 0.0285319f $X=5.895 $Y=1.16 $X2=0 $Y2=0
cc_456 X N_A_814_65#_c_902_n 0.0238338f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_457 N_VGND_c_837_n N_A_814_65#_c_900_n 0.0422287f $X=5.795 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_840_n N_A_814_65#_c_900_n 0.0238173f $X=6 $Y=0 $X2=0 $Y2=0
cc_459 N_VGND_c_831_n N_A_814_65#_c_901_n 0.00500552f $X=3.7 $Y=0.36 $X2=0 $Y2=0
cc_460 N_VGND_c_837_n N_A_814_65#_c_901_n 0.0154127f $X=5.795 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_840_n N_A_814_65#_c_901_n 0.0083587f $X=6 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_c_833_n N_A_814_65#_c_902_n 0.0290385f $X=5.96 $Y=0.47 $X2=0 $Y2=0
cc_463 N_VGND_c_837_n N_A_814_65#_c_902_n 0.0454785f $X=5.795 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_840_n N_A_814_65#_c_902_n 0.0249639f $X=6 $Y=0 $X2=0 $Y2=0
