* File: sky130_fd_sc_lp__or2b_1.pex.spice
* Created: Wed Sep  2 10:29:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2B_1%B_N 3 5 6 7 9 12 13 14 15 20
r41 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.535
+ $Y=0.94 $X2=0.535 $Y2=0.94
r42 15 22 4.82917 $w=4.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.69 $Y=1.665
+ $X2=0.69 $Y2=1.475
r43 14 22 4.48529 $w=4.78e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.295
+ $X2=0.69 $Y2=1.475
r44 14 21 8.846 $w=4.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.69 $Y=1.295
+ $X2=0.69 $Y2=0.94
r45 13 21 0.373774 $w=4.78e-07 $l=1.5e-08 $layer=LI1_cond $X=0.69 $Y=0.925
+ $X2=0.69 $Y2=0.94
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.535 $Y=1.28
+ $X2=0.535 $Y2=0.94
r47 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.28
+ $X2=0.535 $Y2=1.445
r48 10 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.535 $Y=0.925
+ $X2=0.535 $Y2=0.94
r49 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.02 $Y=0.775 $X2=1.02
+ $Y2=0.455
r50 6 10 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.7 $Y=0.85
+ $X2=0.535 $Y2=0.925
r51 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.945 $Y=0.85
+ $X2=1.02 $Y2=0.775
r52 5 6 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.945 $Y=0.85 $X2=0.7
+ $Y2=0.85
r53 3 12 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=0.475 $Y=2.885
+ $X2=0.475 $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_1%A_27_535# 1 2 7 8 9 13 15 17 19 21 24 26 28
+ 30 34 35 37
r81 35 38 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.14 $Y=2.79
+ $X2=0.97 $Y2=2.79
r82 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=2.79 $X2=1.14 $Y2=2.79
r83 32 34 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.14 $Y=2.55 $X2=1.14
+ $Y2=2.79
r84 31 37 2.76166 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.39 $Y=2.465
+ $X2=0.237 $Y2=2.465
r85 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.975 $Y=2.465
+ $X2=1.14 $Y2=2.55
r86 30 31 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.975 $Y=2.465
+ $X2=0.39 $Y2=2.465
r87 26 28 19.2074 $w=3.13e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=0.447
+ $X2=0.805 $Y2=0.447
r88 22 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.237 $Y=2.55
+ $X2=0.237 $Y2=2.465
r89 22 24 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=0.237 $Y=2.55
+ $X2=0.237 $Y2=2.885
r90 21 37 3.70735 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.182 $Y=2.38
+ $X2=0.237 $Y2=2.465
r91 20 26 7.31914 $w=3.15e-07 $l=2.01117e-07 $layer=LI1_cond $X=0.182 $Y=0.605
+ $X2=0.28 $Y2=0.447
r92 20 21 100.956 $w=1.93e-07 $l=1.775e-06 $layer=LI1_cond $X=0.182 $Y=0.605
+ $X2=0.182 $Y2=2.38
r93 15 19 20.4101 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=1.46 $Y=1.725
+ $X2=1.455 $Y2=1.65
r94 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.46 $Y=1.725
+ $X2=1.46 $Y2=2.045
r95 11 19 20.4101 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=1.45 $Y=1.575
+ $X2=1.455 $Y2=1.65
r96 11 13 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.45 $Y=1.575
+ $X2=1.45 $Y2=0.455
r97 10 18 4.07462 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=1.06 $Y=1.65
+ $X2=0.977 $Y2=1.65
r98 9 19 5.30422 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=1.375 $Y=1.65 $X2=1.455
+ $Y2=1.65
r99 9 10 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.375 $Y=1.65
+ $X2=1.06 $Y2=1.65
r100 8 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=2.625
+ $X2=0.97 $Y2=2.79
r101 7 18 56.6087 $w=1.58e-07 $l=1.88467e-07 $layer=POLY_cond $X=0.97 $Y=1.835
+ $X2=0.977 $Y2=1.65
r102 7 8 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.97 $Y=1.835
+ $X2=0.97 $Y2=2.625
r103 2 24 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.885
r104 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.68
+ $Y=0.245 $X2=0.805 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_1%A 4 7 10 11 12 19
c44 11 0 1.97134e-19 $X=1.68 $Y=2.405
r45 16 19 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.68 $Y=2.79
+ $X2=1.82 $Y2=2.79
r46 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=2.79 $X2=1.68 $Y2=2.79
r47 11 12 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=2.405
+ $X2=1.65 $Y2=2.775
r48 9 10 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=1.85 $Y=0.805
+ $X2=1.85 $Y2=0.955
r49 7 9 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.88 $Y=0.455 $X2=1.88
+ $Y2=0.805
r50 4 10 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.82 $Y=2.045
+ $X2=1.82 $Y2=0.955
r51 2 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=2.625
+ $X2=1.82 $Y2=2.79
r52 2 4 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.82 $Y=2.625 $X2=1.82
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_1%A_224_382# 1 2 9 13 16 19 22 23 26 28 30
c57 9 0 1.97134e-19 $X=2.345 $Y=2.465
r58 26 27 16.9324 $w=2.81e-07 $l=3.9e-07 $layer=LI1_cond $X=1.245 $Y=2.045
+ $X2=1.635 $Y2=2.045
r59 23 31 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.292 $Y=1.36
+ $X2=2.292 $Y2=1.525
r60 23 30 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.292 $Y=1.36
+ $X2=2.292 $Y2=1.195
r61 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.27
+ $Y=1.36 $X2=2.27 $Y2=1.36
r62 20 28 0.221902 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.77 $Y=1.36
+ $X2=1.655 $Y2=1.36
r63 20 22 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.77 $Y=1.36 $X2=2.27
+ $Y2=1.36
r64 19 27 3.02819 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=1.88
+ $X2=1.635 $Y2=2.045
r65 18 28 7.38875 $w=2.1e-07 $l=1.74714e-07 $layer=LI1_cond $X=1.635 $Y=1.525
+ $X2=1.655 $Y2=1.36
r66 18 19 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=1.635 $Y=1.525
+ $X2=1.635 $Y2=1.88
r67 14 28 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=1.195
+ $X2=1.655 $Y2=1.36
r68 14 16 37.0786 $w=2.28e-07 $l=7.4e-07 $layer=LI1_cond $X=1.655 $Y=1.195
+ $X2=1.655 $Y2=0.455
r69 13 30 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.405 $Y=0.665
+ $X2=2.405 $Y2=1.195
r70 9 31 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.345 $Y=2.465 $X2=2.345
+ $Y2=1.525
r71 2 26 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.91 $X2=1.245 $Y2=2.045
r72 1 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.525
+ $Y=0.245 $X2=1.665 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_1%VPWR 1 2 9 13 17 19 24 31 32 35 38
r39 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 29 38 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.125 $Y2=3.33
r44 29 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 25 35 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.682 $Y2=3.33
r48 25 27 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 24 38 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.125 $Y2=3.33
r50 24 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 19 35 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.682 $Y2=3.33
r54 19 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r55 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 17 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 13 16 16.1003 $w=3.38e-07 $l=4.75e-07 $layer=LI1_cond $X=2.125 $Y=1.98
+ $X2=2.125 $Y2=2.455
r58 11 38 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=3.33
r59 11 16 26.7774 $w=3.38e-07 $l=7.9e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=2.455
r60 7 35 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.682 $Y=3.245
+ $X2=0.682 $Y2=3.33
r61 7 9 16.9339 $w=2.43e-07 $l=3.6e-07 $layer=LI1_cond $X=0.682 $Y=3.245
+ $X2=0.682 $Y2=2.885
r62 2 16 300 $w=1.7e-07 $l=7.2808e-07 $layer=licon1_PDIFF $count=2 $X=1.895
+ $Y=1.835 $X2=2.13 $Y2=2.455
r63 2 13 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.835 $X2=2.075 $Y2=1.98
r64 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.675 $X2=0.69 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_1%X 1 2 7 8 9 10 11 12 13 24 37
r15 13 44 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.63 $Y=2.775
+ $X2=2.63 $Y2=2.91
r16 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.63 $Y=2.405
+ $X2=2.63 $Y2=2.775
r17 11 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.63 $Y=1.965
+ $X2=2.63 $Y2=1.98
r18 11 47 5.65339 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.63 $Y=1.965
+ $X2=2.63 $Y2=1.815
r19 11 12 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.63 $Y=2.05
+ $X2=2.63 $Y2=2.405
r20 11 37 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=2.63 $Y=2.05 $X2=2.63
+ $Y2=1.98
r21 10 47 6.40246 $w=2.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.66 $Y=1.665
+ $X2=2.66 $Y2=1.815
r22 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=1.295
+ $X2=2.66 $Y2=1.665
r23 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=0.925 $X2=2.66
+ $Y2=1.295
r24 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=0.555 $X2=2.66
+ $Y2=0.925
r25 7 24 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.66 $Y=0.555
+ $X2=2.66 $Y2=0.42
r26 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=2.91
r27 2 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=1.98
r28 1 24 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.48
+ $Y=0.245 $X2=2.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_1%VGND 1 2 9 13 17 19 24 31 32 35 38
r36 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r37 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 29 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.165
+ $Y2=0
r41 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.64
+ $Y2=0
r42 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r43 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r44 25 35 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.255
+ $Y2=0
r45 25 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.68
+ $Y2=0
r46 24 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.165
+ $Y2=0
r47 24 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.68
+ $Y2=0
r48 22 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r49 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 19 35 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=1.255
+ $Y2=0
r51 19 21 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=0.24
+ $Y2=0
r52 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r53 17 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r54 13 15 15.6186 $w=3.78e-07 $l=5.15e-07 $layer=LI1_cond $X=2.165 $Y=0.39
+ $X2=2.165 $Y2=0.905
r55 11 38 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r56 11 13 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.39
r57 7 35 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0
r58 7 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0.455
r59 2 15 182 $w=1.7e-07 $l=7.6857e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.245 $X2=2.19 $Y2=0.905
r60 2 13 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.245 $X2=2.14 $Y2=0.39
r61 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.245 $X2=1.235 $Y2=0.455
.ends

