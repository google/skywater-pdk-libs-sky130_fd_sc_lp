* File: sky130_fd_sc_lp__o2bb2ai_2.spice
* Created: Fri Aug 28 11:12:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2ai_2.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2ai_2  VNB VPB A1_N A2_N B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A1_N_M1015_g N_A_125_69#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1008 N_A_125_69#_M1015_s N_A2_N_M1008_g N_A_125_367#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1018 N_A_125_69#_M1018_d N_A2_N_M1018_g N_A_125_367#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_A1_N_M1017_g N_A_125_69#_M1018_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A_125_367#_M1000_g N_A_502_69#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1006 N_Y_M1000_d N_A_125_367#_M1006_g N_A_502_69#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=5.712 M=1 R=5.6 SA=75000.6
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_B1_M1012_g N_A_502_69#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=5.712 M=1 R=5.6 SA=75001.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1003 N_A_502_69#_M1003_d N_B2_M1003_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1010 N_A_502_69#_M1003_d N_B2_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1010_s N_B1_M1016_g N_A_502_69#_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_A1_N_M1001_g N_A_125_367#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1009 N_A_125_367#_M1001_s N_A2_N_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1014 N_A_125_367#_M1014_d N_A2_N_M1014_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_N_M1007_g N_A_125_367#_M1014_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.5418 AS=0.1764 PD=2.12 PS=1.54 NRD=68.0044 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75003.4 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_A_125_367#_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.5418 PD=1.54 PS=2.12 NRD=0 NRS=22.655 M=1 R=8.4 SA=75002.5
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1004_d N_A_125_367#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75002.9
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1019_s N_B1_M1011_g N_A_765_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75003.4 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1002 N_A_765_367#_M1011_s N_B2_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75003.8
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_A_765_367#_M1005_d N_B2_M1005_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75004.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_B1_M1013_g N_A_765_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__o2bb2ai_2.pxi.spice"
*
.ends
*
*
