* File: sky130_fd_sc_lp__invlp_1.spice
* Created: Fri Aug 28 10:39:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__invlp_1.pex.spice"
.subckt sky130_fd_sc_lp__invlp_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 A_124_47# N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2394 PD=1.08 PS=2.25 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g A_124_47# VNB NSHORT L=0.15 W=0.84 AD=0.2394
+ AS=0.1008 PD=2.25 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1000 A_130_367# N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.3591 PD=1.47 PS=3.09 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_130_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.3591
+ AS=0.1323 PD=3.09 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__invlp_1.pxi.spice"
*
.ends
*
*
