* File: sky130_fd_sc_lp__a221oi_1.pex.spice
* Created: Fri Aug 28 09:53:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221OI_1%C1 3 7 9 10 17
r33 15 17 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.64 $Y=1.375 $X2=0.71
+ $Y2=1.375
r34 13 15 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.375
+ $X2=0.64 $Y2=1.375
r35 9 10 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.702 $Y=1.295
+ $X2=0.702 $Y2=1.665
r36 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.375 $X2=0.71 $Y2=1.375
r37 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.21
+ $X2=0.64 $Y2=1.375
r38 5 7 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.64 $Y=1.21 $X2=0.64
+ $Y2=0.655
r39 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=1.375
r40 1 3 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%B2 3 6 8 11 12 13
r37 11 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.32 $Y=1.35
+ $X2=1.32 $Y2=1.515
r38 11 13 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.32 $Y=1.35
+ $X2=1.32 $Y2=1.185
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.305
+ $Y=1.35 $X2=1.305 $Y2=1.35
r40 8 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.35
+ $X2=1.305 $Y2=1.35
r41 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.425 $Y=2.465
+ $X2=1.425 $Y2=1.515
r42 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.425 $Y=0.655
+ $X2=1.425 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%B1 3 6 8 11 12 13
r32 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.35
+ $X2=1.875 $Y2=1.185
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.875
+ $Y=1.35 $X2=1.875 $Y2=1.35
r34 8 12 7.36808 $w=3.03e-07 $l=1.95e-07 $layer=LI1_cond $X=1.68 $Y=1.362
+ $X2=1.875 $Y2=1.362
r35 4 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.515
+ $X2=1.875 $Y2=1.35
r36 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.875 $Y=1.515
+ $X2=1.875 $Y2=2.465
r37 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.785 $Y=0.655
+ $X2=1.785 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%A1 3 6 8 9 10 15 17
r32 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.515
r33 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.185
r34 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.35 $X2=2.415 $Y2=1.35
r35 10 16 1.4914 $w=4.23e-07 $l=5.5e-08 $layer=LI1_cond $X=2.522 $Y=1.295
+ $X2=2.522 $Y2=1.35
r36 10 26 4.23752 $w=4.23e-07 $l=1.1e-07 $layer=LI1_cond $X=2.522 $Y=1.295
+ $X2=2.522 $Y2=1.185
r37 9 26 10.5135 $w=2.83e-07 $l=2.6e-07 $layer=LI1_cond $X=2.592 $Y=0.925
+ $X2=2.592 $Y2=1.185
r38 8 9 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.592 $Y=0.555
+ $X2=2.592 $Y2=0.925
r39 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.355 $Y=2.465
+ $X2=2.355 $Y2=1.515
r40 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.325 $Y=0.655
+ $X2=2.325 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%A2 3 6 8 11 13
r23 11 14 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.972 $Y=1.35
+ $X2=2.972 $Y2=1.515
r24 11 13 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.972 $Y=1.35
+ $X2=2.972 $Y2=1.185
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.35 $X2=2.99 $Y2=1.35
r26 8 12 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.35 $X2=2.99
+ $Y2=1.35
r27 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.865 $Y=2.465
+ $X2=2.865 $Y2=1.515
r28 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.865 $Y=0.655
+ $X2=2.865 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%Y 1 2 3 10 14 16 17 18 19 20 21 22 33
r32 22 51 5.45894 $w=2.83e-07 $l=1.35e-07 $layer=LI1_cond $X=0.232 $Y=2.775
+ $X2=0.232 $Y2=2.91
r33 21 22 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.232 $Y=2.405
+ $X2=0.232 $Y2=2.775
r34 20 21 17.1856 $w=2.83e-07 $l=4.25e-07 $layer=LI1_cond $X=0.232 $Y=1.98
+ $X2=0.232 $Y2=2.405
r35 19 20 12.7375 $w=2.83e-07 $l=3.15e-07 $layer=LI1_cond $X=0.232 $Y=1.665
+ $X2=0.232 $Y2=1.98
r36 18 19 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.232 $Y=1.295
+ $X2=0.232 $Y2=1.665
r37 18 38 11.3222 $w=2.83e-07 $l=2.8e-07 $layer=LI1_cond $X=0.232 $Y=1.295
+ $X2=0.232 $Y2=1.015
r38 17 31 2.68319 $w=3.57e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=0.93
+ $X2=0.305 $Y2=0.845
r39 17 38 2.68319 $w=3.57e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.305 $Y=0.93
+ $X2=0.232 $Y2=1.015
r40 17 31 0.080403 $w=4.28e-07 $l=3e-09 $layer=LI1_cond $X=0.305 $Y=0.842
+ $X2=0.305 $Y2=0.845
r41 16 17 7.69189 $w=4.28e-07 $l=2.87e-07 $layer=LI1_cond $X=0.305 $Y=0.555
+ $X2=0.305 $Y2=0.842
r42 16 33 3.35013 $w=4.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.305 $Y=0.555
+ $X2=0.305 $Y2=0.43
r43 12 14 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.055 $Y=0.845
+ $X2=2.055 $Y2=0.38
r44 11 17 4.11427 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.52 $Y=0.93
+ $X2=0.305 $Y2=0.93
r45 10 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.89 $Y=0.93
+ $X2=2.055 $Y2=0.845
r46 10 11 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.89 $Y=0.93
+ $X2=0.52 $Y2=0.93
r47 3 51 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r48 3 20 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r49 2 14 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.235 $X2=2.055 $Y2=0.38
r50 1 33 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=0.3 $Y=0.235
+ $X2=0.425 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%A_110_367# 1 2 7 9 11 15
r20 15 18 33.8377 $w=2.33e-07 $l=6.9e-07 $layer=LI1_cond $X=1.662 $Y=2.21
+ $X2=1.662 $Y2=2.9
r21 13 18 0.245201 $w=2.33e-07 $l=5e-09 $layer=LI1_cond $X=1.662 $Y=2.905
+ $X2=1.662 $Y2=2.9
r22 12 20 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.855 $Y=2.99
+ $X2=0.7 $Y2=2.99
r23 11 13 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=1.545 $Y=2.99
+ $X2=1.662 $Y2=2.905
r24 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.545 $Y=2.99
+ $X2=0.855 $Y2=2.99
r25 7 20 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.905 $X2=0.7
+ $Y2=2.99
r26 7 9 30.484 $w=3.08e-07 $l=8.2e-07 $layer=LI1_cond $X=0.7 $Y=2.905 $X2=0.7
+ $Y2=2.085
r27 2 18 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.9
r28 2 15 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.21
r29 1 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.91
r30 1 9 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%A_217_367# 1 2 3 12 14 15 18 22 26 30
r44 26 28 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.11 $Y=1.98
+ $X2=3.11 $Y2=2.91
r45 24 26 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.11 $Y=1.875
+ $X2=3.11 $Y2=1.98
r46 23 30 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.27 $Y=1.79 $X2=2.11
+ $Y2=1.79
r47 22 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.975 $Y=1.79
+ $X2=3.11 $Y2=1.875
r48 22 23 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.975 $Y=1.79
+ $X2=2.27 $Y2=1.79
r49 18 20 33.4929 $w=3.18e-07 $l=9.3e-07 $layer=LI1_cond $X=2.11 $Y=1.98
+ $X2=2.11 $Y2=2.91
r50 16 30 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=1.875
+ $X2=2.11 $Y2=1.79
r51 16 18 3.78145 $w=3.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.11 $Y=1.875
+ $X2=2.11 $Y2=1.98
r52 14 30 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.95 $Y=1.79 $X2=2.11
+ $Y2=1.79
r53 14 15 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.95 $Y=1.79
+ $X2=1.375 $Y2=1.79
r54 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.21 $Y=1.875
+ $X2=1.375 $Y2=1.79
r55 10 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.21 $Y=1.875
+ $X2=1.21 $Y2=1.98
r56 3 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=2.91
r57 3 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=1.98
r58 2 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.09 $Y2=2.91
r59 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.09 $Y2=1.98
r60 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%VPWR 1 6 10 12 22 23 26
r36 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 23 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 20 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.605 $Y2=3.33
r40 20 22 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 19 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 12 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=3.33
+ $X2=2.605 $Y2=3.33
r46 12 18 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 10 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 6 9 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=2.605 $Y=2.13
+ $X2=2.605 $Y2=2.95
r50 4 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=3.245
+ $X2=2.605 $Y2=3.33
r51 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.605 $Y=3.245
+ $X2=2.605 $Y2=2.95
r52 1 9 400 $w=1.7e-07 $l=1.19931e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.835 $X2=2.605 $Y2=2.95
r53 1 6 400 $w=1.7e-07 $l=3.72357e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.835 $X2=2.605 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_1%VGND 1 2 7 9 11 13 15 34
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r35 26 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r36 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r37 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 18 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r39 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r40 15 33 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r41 15 21 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r42 13 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r43 13 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r44 13 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 9 33 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r46 9 11 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.38
r47 7 30 9.60355 $w=6.83e-07 $l=5.5e-07 $layer=LI1_cond $X=1.032 $Y=0 $X2=1.032
+ $Y2=0.55
r48 7 16 9.17904 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=1.032 $Y=0 $X2=1.375
+ $Y2=0
r49 7 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 7 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.38
r52 1 30 91 $w=1.7e-07 $l=6.33206e-07 $layer=licon1_NDIFF $count=2 $X=0.715
+ $Y=0.235 $X2=1.21 $Y2=0.55
.ends

