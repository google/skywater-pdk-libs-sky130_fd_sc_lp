* File: sky130_fd_sc_lp__sdfbbp_1.pxi.spice
* Created: Fri Aug 28 11:27:30 2020
* 
x_PM_SKY130_FD_SC_LP__SDFBBP_1%SCD N_SCD_M1037_g N_SCD_M1033_g N_SCD_c_350_n
+ N_SCD_c_354_n N_SCD_c_355_n N_SCD_c_356_n SCD N_SCD_c_351_n N_SCD_c_352_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%SCD
x_PM_SKY130_FD_SC_LP__SDFBBP_1%D N_D_M1019_g N_D_M1005_g D N_D_c_392_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%D
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_332_93# N_A_332_93#_M1034_d N_A_332_93#_M1038_d
+ N_A_332_93#_c_433_n N_A_332_93#_M1003_g N_A_332_93#_M1041_g
+ N_A_332_93#_c_434_n N_A_332_93#_c_435_n N_A_332_93#_c_436_n
+ N_A_332_93#_c_442_n N_A_332_93#_c_443_n N_A_332_93#_c_437_n
+ N_A_332_93#_c_438_n N_A_332_93#_c_445_n N_A_332_93#_c_446_n
+ N_A_332_93#_c_439_n N_A_332_93#_c_440_n N_A_332_93#_c_449_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_332_93#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%SCE N_SCE_M1013_g N_SCE_M1032_g N_SCE_c_525_n
+ N_SCE_c_526_n N_SCE_M1034_g N_SCE_c_528_n N_SCE_c_529_n N_SCE_M1038_g
+ N_SCE_c_535_n N_SCE_c_536_n N_SCE_c_530_n N_SCE_c_538_n SCE N_SCE_c_532_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%SCE
x_PM_SKY130_FD_SC_LP__SDFBBP_1%CLK N_CLK_M1015_g N_CLK_M1006_g N_CLK_c_625_n
+ N_CLK_c_626_n CLK CLK N_CLK_c_623_n PM_SKY130_FD_SC_LP__SDFBBP_1%CLK
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_893_101# N_A_893_101#_M1022_s
+ N_A_893_101#_M1042_s N_A_893_101#_c_663_n N_A_893_101#_c_664_n
+ N_A_893_101#_c_665_n N_A_893_101#_M1012_g N_A_893_101#_c_667_n
+ N_A_893_101#_c_668_n N_A_893_101#_M1023_g N_A_893_101#_c_681_n
+ N_A_893_101#_M1029_g N_A_893_101#_M1018_g N_A_893_101#_c_671_n
+ N_A_893_101#_c_672_n N_A_893_101#_c_683_n N_A_893_101#_c_684_n
+ N_A_893_101#_c_685_n N_A_893_101#_c_686_n N_A_893_101#_c_673_n
+ N_A_893_101#_c_674_n N_A_893_101#_c_675_n N_A_893_101#_c_676_n
+ N_A_893_101#_c_677_n N_A_893_101#_c_678_n N_A_893_101#_c_679_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_893_101#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_1297_290# N_A_1297_290#_M1001_d
+ N_A_1297_290#_M1040_d N_A_1297_290#_M1016_g N_A_1297_290#_M1010_g
+ N_A_1297_290#_M1031_g N_A_1297_290#_c_839_n N_A_1297_290#_c_840_n
+ N_A_1297_290#_M1008_g N_A_1297_290#_c_851_n N_A_1297_290#_c_852_n
+ N_A_1297_290#_c_972_p N_A_1297_290#_c_866_n N_A_1297_290#_c_887_p
+ N_A_1297_290#_c_867_n N_A_1297_290#_c_842_n N_A_1297_290#_c_854_n
+ N_A_1297_290#_c_843_n N_A_1297_290#_c_844_n N_A_1297_290#_c_845_n
+ N_A_1297_290#_c_880_n N_A_1297_290#_c_903_p N_A_1297_290#_c_846_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_1297_290#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%SET_B N_SET_B_M1026_g N_SET_B_M1040_g
+ N_SET_B_M1011_g N_SET_B_c_1019_n N_SET_B_M1020_g N_SET_B_c_1027_n SET_B
+ N_SET_B_c_1029_n N_SET_B_c_1030_n N_SET_B_c_1021_n N_SET_B_c_1022_n
+ N_SET_B_c_1033_n N_SET_B_c_1034_n PM_SKY130_FD_SC_LP__SDFBBP_1%SET_B
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_1216_457# N_A_1216_457#_M1004_d
+ N_A_1216_457#_M1012_d N_A_1216_457#_M1001_g N_A_1216_457#_M1024_g
+ N_A_1216_457#_c_1154_n N_A_1216_457#_c_1155_n N_A_1216_457#_c_1156_n
+ N_A_1216_457#_c_1157_n N_A_1216_457#_c_1158_n N_A_1216_457#_c_1159_n
+ N_A_1216_457#_c_1160_n N_A_1216_457#_c_1161_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_1216_457#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_1650_21# N_A_1650_21#_M1002_s
+ N_A_1650_21#_M1000_s N_A_1650_21#_c_1248_n N_A_1650_21#_M1007_g
+ N_A_1650_21#_M1046_g N_A_1650_21#_M1014_g N_A_1650_21#_c_1251_n
+ N_A_1650_21#_M1047_g N_A_1650_21#_c_1252_n N_A_1650_21#_c_1253_n
+ N_A_1650_21#_c_1254_n N_A_1650_21#_c_1255_n N_A_1650_21#_c_1256_n
+ N_A_1650_21#_c_1406_p N_A_1650_21#_c_1257_n N_A_1650_21#_c_1258_n
+ N_A_1650_21#_c_1259_n N_A_1650_21#_c_1260_n N_A_1650_21#_c_1261_n
+ N_A_1650_21#_c_1262_n N_A_1650_21#_c_1263_n N_A_1650_21#_c_1264_n
+ N_A_1650_21#_c_1265_n N_A_1650_21#_c_1266_n N_A_1650_21#_c_1267_n
+ N_A_1650_21#_c_1268_n PM_SKY130_FD_SC_LP__SDFBBP_1%A_1650_21#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_755_106# N_A_755_106#_M1015_d
+ N_A_755_106#_M1006_d N_A_755_106#_c_1421_n N_A_755_106#_c_1422_n
+ N_A_755_106#_c_1423_n N_A_755_106#_M1022_g N_A_755_106#_M1042_g
+ N_A_755_106#_c_1425_n N_A_755_106#_c_1436_n N_A_755_106#_c_1437_n
+ N_A_755_106#_c_1426_n N_A_755_106#_c_1427_n N_A_755_106#_c_1428_n
+ N_A_755_106#_c_1429_n N_A_755_106#_M1004_g N_A_755_106#_M1043_g
+ N_A_755_106#_c_1439_n N_A_755_106#_M1035_g N_A_755_106#_c_1441_n
+ N_A_755_106#_c_1442_n N_A_755_106#_M1027_g N_A_755_106#_c_1431_n
+ N_A_755_106#_c_1444_n N_A_755_106#_c_1432_n N_A_755_106#_c_1433_n
+ N_A_755_106#_c_1446_n N_A_755_106#_c_1434_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_755_106#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_2064_453# N_A_2064_453#_M1028_d
+ N_A_2064_453#_M1020_d N_A_2064_453#_M1017_g N_A_2064_453#_M1009_g
+ N_A_2064_453#_M1036_g N_A_2064_453#_M1045_g N_A_2064_453#_c_1583_n
+ N_A_2064_453#_M1039_g N_A_2064_453#_M1025_g N_A_2064_453#_c_1596_n
+ N_A_2064_453#_c_1586_n N_A_2064_453#_c_1597_n N_A_2064_453#_c_1598_n
+ N_A_2064_453#_c_1599_n N_A_2064_453#_c_1600_n N_A_2064_453#_c_1648_p
+ N_A_2064_453#_c_1587_n N_A_2064_453#_c_1602_n N_A_2064_453#_c_1588_n
+ N_A_2064_453#_c_1638_n N_A_2064_453#_c_1589_n N_A_2064_453#_c_1642_n
+ N_A_2064_453#_c_1590_n N_A_2064_453#_c_1591_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_2064_453#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_1861_431# N_A_1861_431#_M1018_d
+ N_A_1861_431#_M1035_d N_A_1861_431#_M1028_g N_A_1861_431#_M1021_g
+ N_A_1861_431#_c_1765_n N_A_1861_431#_c_1754_n N_A_1861_431#_c_1755_n
+ N_A_1861_431#_c_1756_n N_A_1861_431#_c_1757_n N_A_1861_431#_c_1758_n
+ N_A_1861_431#_c_1764_n N_A_1861_431#_c_1759_n N_A_1861_431#_c_1760_n
+ N_A_1861_431#_c_1761_n PM_SKY130_FD_SC_LP__SDFBBP_1%A_1861_431#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%RESET_B N_RESET_B_M1002_g N_RESET_B_M1000_g
+ RESET_B N_RESET_B_c_1875_n N_RESET_B_c_1876_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%RESET_B
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_2892_137# N_A_2892_137#_M1039_s
+ N_A_2892_137#_M1025_s N_A_2892_137#_M1030_g N_A_2892_137#_M1044_g
+ N_A_2892_137#_c_1910_n N_A_2892_137#_c_1915_n N_A_2892_137#_c_1911_n
+ N_A_2892_137#_c_1912_n N_A_2892_137#_c_1913_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_2892_137#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_27_481# N_A_27_481#_M1037_s N_A_27_481#_M1041_d
+ N_A_27_481#_c_1960_n N_A_27_481#_c_1961_n N_A_27_481#_c_1962_n
+ N_A_27_481#_c_1963_n N_A_27_481#_c_1964_n N_A_27_481#_c_1965_n
+ N_A_27_481#_c_1966_n PM_SKY130_FD_SC_LP__SDFBBP_1%A_27_481#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%VPWR N_VPWR_M1037_d N_VPWR_M1038_s N_VPWR_M1006_s
+ N_VPWR_M1042_d N_VPWR_M1016_d N_VPWR_M1046_d N_VPWR_M1017_d N_VPWR_M1014_d
+ N_VPWR_M1000_d N_VPWR_M1025_d N_VPWR_c_2011_n N_VPWR_c_2012_n N_VPWR_c_2013_n
+ N_VPWR_c_2014_n N_VPWR_c_2015_n N_VPWR_c_2016_n N_VPWR_c_2017_n
+ N_VPWR_c_2018_n N_VPWR_c_2019_n N_VPWR_c_2020_n N_VPWR_c_2021_n
+ N_VPWR_c_2022_n N_VPWR_c_2023_n N_VPWR_c_2024_n N_VPWR_c_2025_n
+ N_VPWR_c_2026_n N_VPWR_c_2027_n VPWR N_VPWR_c_2028_n N_VPWR_c_2029_n
+ N_VPWR_c_2030_n N_VPWR_c_2031_n N_VPWR_c_2032_n N_VPWR_c_2033_n
+ N_VPWR_c_2034_n N_VPWR_c_2010_n N_VPWR_c_2036_n N_VPWR_c_2037_n
+ N_VPWR_c_2038_n N_VPWR_c_2039_n N_VPWR_c_2040_n N_VPWR_c_2041_n
+ N_VPWR_c_2042_n PM_SKY130_FD_SC_LP__SDFBBP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_204_119# N_A_204_119#_M1013_d
+ N_A_204_119#_M1004_s N_A_204_119#_M1005_d N_A_204_119#_M1012_s
+ N_A_204_119#_c_2199_n N_A_204_119#_c_2200_n N_A_204_119#_c_2201_n
+ N_A_204_119#_c_2218_n N_A_204_119#_c_2202_n N_A_204_119#_c_2203_n
+ N_A_204_119#_c_2204_n N_A_204_119#_c_2205_n N_A_204_119#_c_2206_n
+ N_A_204_119#_c_2207_n N_A_204_119#_c_2208_n N_A_204_119#_c_2209_n
+ N_A_204_119#_c_2210_n N_A_204_119#_c_2211_n N_A_204_119#_c_2326_n
+ N_A_204_119#_c_2212_n N_A_204_119#_c_2213_n N_A_204_119#_c_2214_n
+ N_A_204_119#_c_2220_n N_A_204_119#_c_2215_n N_A_204_119#_c_2221_n
+ N_A_204_119#_c_2216_n N_A_204_119#_c_2217_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%A_204_119#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%Q_N N_Q_N_M1036_d N_Q_N_M1045_d N_Q_N_c_2395_n
+ N_Q_N_c_2396_n N_Q_N_c_2398_n N_Q_N_c_2397_n Q_N Q_N Q_N
+ PM_SKY130_FD_SC_LP__SDFBBP_1%Q_N
x_PM_SKY130_FD_SC_LP__SDFBBP_1%Q N_Q_M1030_d N_Q_M1044_d N_Q_c_2432_n
+ N_Q_c_2433_n N_Q_c_2429_n Q Q N_Q_c_2431_n Q PM_SKY130_FD_SC_LP__SDFBBP_1%Q
x_PM_SKY130_FD_SC_LP__SDFBBP_1%VGND N_VGND_M1033_s N_VGND_M1003_d N_VGND_M1015_s
+ N_VGND_M1022_d N_VGND_M1010_d N_VGND_M1008_s N_VGND_M1009_d N_VGND_M1002_d
+ N_VGND_M1039_d N_VGND_c_2454_n N_VGND_c_2455_n N_VGND_c_2456_n N_VGND_c_2457_n
+ N_VGND_c_2458_n N_VGND_c_2459_n N_VGND_c_2460_n N_VGND_c_2461_n
+ N_VGND_c_2462_n N_VGND_c_2463_n N_VGND_c_2464_n N_VGND_c_2465_n
+ N_VGND_c_2466_n N_VGND_c_2467_n N_VGND_c_2468_n N_VGND_c_2469_n
+ N_VGND_c_2470_n N_VGND_c_2471_n N_VGND_c_2472_n N_VGND_c_2473_n
+ N_VGND_c_2474_n N_VGND_c_2475_n N_VGND_c_2476_n N_VGND_c_2477_n VGND
+ N_VGND_c_2478_n N_VGND_c_2479_n N_VGND_c_2480_n N_VGND_c_2481_n
+ PM_SKY130_FD_SC_LP__SDFBBP_1%VGND
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_1492_47# N_A_1492_47#_M1026_d
+ N_A_1492_47#_M1007_d N_A_1492_47#_c_2640_n N_A_1492_47#_c_2646_n
+ N_A_1492_47#_c_2639_n PM_SKY130_FD_SC_LP__SDFBBP_1%A_1492_47#
x_PM_SKY130_FD_SC_LP__SDFBBP_1%A_2279_57# N_A_2279_57#_M1011_d
+ N_A_2279_57#_M1047_d N_A_2279_57#_c_2669_n N_A_2279_57#_c_2670_n
+ N_A_2279_57#_c_2671_n PM_SKY130_FD_SC_LP__SDFBBP_1%A_2279_57#
cc_1 VNB N_SCD_M1033_g 0.0237224f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.805
cc_2 VNB N_SCD_c_350_n 0.025908f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.31
cc_3 VNB N_SCD_c_351_n 0.0264991f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_4 VNB N_SCD_c_352_n 0.0228759f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_5 VNB N_D_M1019_g 0.0361293f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.27
cc_6 VNB D 8.42075e-19 $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.805
cc_7 VNB N_D_c_392_n 0.0180689f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.885
cc_8 VNB N_A_332_93#_c_433_n 0.01373f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.16
cc_9 VNB N_A_332_93#_c_434_n 0.0240935f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.72
cc_10 VNB N_A_332_93#_c_435_n 0.00679722f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.885
cc_11 VNB N_A_332_93#_c_436_n 0.0163353f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.27
cc_12 VNB N_A_332_93#_c_437_n 0.00337939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_332_93#_c_438_n 0.00599536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_332_93#_c_439_n 0.00391378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_332_93#_c_440_n 0.0176634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_M1013_g 0.0520831f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.725
cc_17 VNB N_SCE_c_525_n 0.113452f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.31
cc_18 VNB N_SCE_c_526_n 0.0125534f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.16
cc_19 VNB N_SCE_M1034_g 0.0278666f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.12
cc_20 VNB N_SCE_c_528_n 0.0364944f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.27
cc_21 VNB N_SCE_c_529_n 0.00674785f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_SCE_c_530_n 0.0256362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB SCE 0.00330031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_532_n 0.0132779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_CLK_M1015_g 0.045168f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.27
cc_26 VNB CLK 0.0017134f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.12
cc_27 VNB N_CLK_c_623_n 0.0170143f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_28 VNB N_A_893_101#_c_663_n 0.0197239f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.16
cc_29 VNB N_A_893_101#_c_664_n 0.010809f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.805
cc_30 VNB N_A_893_101#_c_665_n 0.012337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_893_101#_M1012_g 0.00493202f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.31
cc_32 VNB N_A_893_101#_c_667_n 0.0349516f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.885
cc_33 VNB N_A_893_101#_c_668_n 0.00766443f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.12
cc_34 VNB N_A_893_101#_M1023_g 0.031299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_893_101#_M1018_g 0.0246343f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.55
cc_36 VNB N_A_893_101#_c_671_n 0.00621012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_893_101#_c_672_n 0.00907068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_893_101#_c_673_n 0.0479146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_893_101#_c_674_n 0.00201427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_893_101#_c_675_n 0.00225379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_893_101#_c_676_n 0.00562986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_893_101#_c_677_n 0.0081646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_893_101#_c_678_n 0.0288737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_893_101#_c_679_n 0.00812646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1297_290#_M1010_g 0.0529826f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.31
cc_46 VNB N_A_1297_290#_c_839_n 0.00863259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1297_290#_c_840_n 0.00734103f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.38
cc_48 VNB N_A_1297_290#_M1008_g 0.0244232f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.55
cc_49 VNB N_A_1297_290#_c_842_n 0.00504284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1297_290#_c_843_n 0.00423977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1297_290#_c_844_n 0.0459136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1297_290#_c_845_n 0.00142916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1297_290#_c_846_n 0.0257453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SET_B_M1026_g 0.0356184f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.27
cc_55 VNB N_SET_B_M1011_g 0.0570495f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.31
cc_56 VNB N_SET_B_c_1019_n 0.0114519f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.31
cc_57 VNB SET_B 0.00521344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_1021_n 3.26246e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SET_B_c_1022_n 0.0200469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1216_457#_M1001_g 0.0196278f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=0.805
cc_61 VNB N_A_1216_457#_c_1154_n 0.0216853f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.27
cc_62 VNB N_A_1216_457#_c_1155_n 0.00857204f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_63 VNB N_A_1216_457#_c_1156_n 0.00102975f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.38
cc_64 VNB N_A_1216_457#_c_1157_n 0.00755367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1216_457#_c_1158_n 0.0212599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1216_457#_c_1159_n 4.736e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1216_457#_c_1160_n 0.0016899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1216_457#_c_1161_n 0.01554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1650_21#_c_1248_n 0.0196094f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.16
cc_70 VNB N_A_1650_21#_M1046_g 0.0174364f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.16
cc_71 VNB N_A_1650_21#_M1014_g 0.0079019f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.12
cc_72 VNB N_A_1650_21#_c_1251_n 0.0659823f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_73 VNB N_A_1650_21#_c_1252_n 0.0389216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1650_21#_c_1253_n 0.00342877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1650_21#_c_1254_n 0.0522875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1650_21#_c_1255_n 0.00752928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1650_21#_c_1256_n 0.00292959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1650_21#_c_1257_n 0.0133459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1650_21#_c_1258_n 0.00140658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1650_21#_c_1259_n 0.00109883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1650_21#_c_1260_n 0.0197185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1650_21#_c_1261_n 0.0018134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1650_21#_c_1262_n 0.0039793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1650_21#_c_1263_n 0.00119558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1650_21#_c_1264_n 0.00297235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1650_21#_c_1265_n 0.00916654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1650_21#_c_1266_n 0.00186502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1650_21#_c_1267_n 0.00222592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1650_21#_c_1268_n 0.00318053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_755_106#_c_1421_n 0.0304256f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.16
cc_91 VNB N_A_755_106#_c_1422_n 0.016379f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.805
cc_92 VNB N_A_755_106#_c_1423_n 0.0210781f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=0.805
cc_93 VNB N_A_755_106#_M1042_g 0.0278313f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.885
cc_94 VNB N_A_755_106#_c_1425_n 0.0369398f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.12
cc_95 VNB N_A_755_106#_c_1426_n 0.00958557f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.38
cc_96 VNB N_A_755_106#_c_1427_n 0.0279341f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_97 VNB N_A_755_106#_c_1428_n 0.0115669f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.55
cc_98 VNB N_A_755_106#_c_1429_n 0.0170876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_755_106#_M1027_g 0.0453628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_755_106#_c_1431_n 0.00382064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_755_106#_c_1432_n 0.00991534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_755_106#_c_1433_n 0.0339048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_755_106#_c_1434_n 7.31569e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2064_453#_M1009_g 0.0507937f $X=-0.19 $Y=-0.245 $X2=0.425
+ $Y2=1.31
cc_105 VNB N_A_2064_453#_M1036_g 0.0272416f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.27
cc_106 VNB N_A_2064_453#_M1045_g 0.0010556f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.38
cc_107 VNB N_A_2064_453#_c_1583_n 0.0597441f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.55
cc_108 VNB N_A_2064_453#_M1039_g 0.0231097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2064_453#_M1025_g 0.0138328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2064_453#_c_1586_n 0.00454738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2064_453#_c_1587_n 0.0065316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2064_453#_c_1588_n 2.66907e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2064_453#_c_1589_n 0.010744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2064_453#_c_1590_n 0.00451298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2064_453#_c_1591_n 0.0317134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1861_431#_M1028_g 0.0564116f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=0.805
cc_117 VNB N_A_1861_431#_M1021_g 0.00163545f $X=-0.19 $Y=-0.245 $X2=0.425
+ $Y2=1.31
cc_118 VNB N_A_1861_431#_c_1754_n 0.00668176f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.27
cc_119 VNB N_A_1861_431#_c_1755_n 0.00311378f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.38
cc_120 VNB N_A_1861_431#_c_1756_n 0.0012905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_1861_431#_c_1757_n 0.0246853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_1861_431#_c_1758_n 0.00213506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_1861_431#_c_1759_n 0.00408108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1861_431#_c_1760_n 0.00330243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_1861_431#_c_1761_n 0.0355384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_RESET_B_M1000_g 0.00522925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB RESET_B 0.00364319f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.805
cc_128 VNB N_RESET_B_c_1875_n 0.0346985f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.31
cc_129 VNB N_RESET_B_c_1876_n 0.020579f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.31
cc_130 VNB N_A_2892_137#_M1030_g 0.0292364f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=0.805
cc_131 VNB N_A_2892_137#_M1044_g 0.00114499f $X=-0.19 $Y=-0.245 $X2=0.425
+ $Y2=1.31
cc_132 VNB N_A_2892_137#_c_1910_n 0.0044825f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.27
cc_133 VNB N_A_2892_137#_c_1911_n 0.00708653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_2892_137#_c_1912_n 0.0345037f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.55
cc_135 VNB N_A_2892_137#_c_1913_n 0.00192268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VPWR_c_2010_n 0.661241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_204_119#_c_2199_n 0.00264581f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.885
cc_138 VNB N_A_204_119#_c_2200_n 0.0155507f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.27
cc_139 VNB N_A_204_119#_c_2201_n 0.00303081f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_140 VNB N_A_204_119#_c_2202_n 0.00319941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_204_119#_c_2203_n 0.00313518f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.55
cc_142 VNB N_A_204_119#_c_2204_n 0.0129702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_204_119#_c_2205_n 0.00254967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_204_119#_c_2206_n 0.0136022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_204_119#_c_2207_n 0.0285264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_A_204_119#_c_2208_n 5.11203e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_204_119#_c_2209_n 0.00787625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_A_204_119#_c_2210_n 0.0273987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_204_119#_c_2211_n 0.00288738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_A_204_119#_c_2212_n 0.00484514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_A_204_119#_c_2213_n 0.00110246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_A_204_119#_c_2214_n 0.00595509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_204_119#_c_2215_n 0.0055886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_204_119#_c_2216_n 0.00556684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_A_204_119#_c_2217_n 0.00126889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_Q_N_c_2395_n 0.0111865f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.805
cc_157 VNB N_Q_N_c_2396_n 0.00555276f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.31
cc_158 VNB N_Q_N_c_2397_n 0.00548581f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.27
cc_159 VNB N_Q_c_2429_n 0.0251675f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.885
cc_160 VNB Q 0.0137223f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.27
cc_161 VNB N_Q_c_2431_n 0.0290706f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.55
cc_162 VNB N_VGND_c_2454_n 0.0141307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2455_n 0.0424769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2456_n 0.01063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2457_n 0.0147907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2458_n 0.0116278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2459_n 0.00713304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2460_n 0.00811363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2461_n 0.00962116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2462_n 0.016851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2463_n 0.0153251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2464_n 0.0379769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2465_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2466_n 0.0300138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2467_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2468_n 0.0437247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2469_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2470_n 0.04331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2471_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2472_n 0.0416977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2473_n 0.00552821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2474_n 0.0388274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2475_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2476_n 0.0346791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2477_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2478_n 0.0589651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2479_n 0.0191143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2480_n 0.82215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_VGND_c_2481_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_A_1492_47#_c_2639_n 0.00210877f $X=-0.19 $Y=-0.245 $X2=0.425
+ $Y2=1.16
cc_191 VNB N_A_2279_57#_c_2669_n 0.00332359f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=1.16
cc_192 VNB N_A_2279_57#_c_2670_n 0.00205429f $X=-0.19 $Y=-0.245 $X2=0.555
+ $Y2=0.805
cc_193 VNB N_A_2279_57#_c_2671_n 0.00239641f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.72
cc_194 VPB N_SCD_M1037_g 0.0233016f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.725
cc_195 VPB N_SCD_c_354_n 0.0168207f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.885
cc_196 VPB N_SCD_c_355_n 0.0187564f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.12
cc_197 VPB N_SCD_c_356_n 0.0108221f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.27
cc_198 VPB N_SCD_c_351_n 0.00472232f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_199 VPB N_SCD_c_352_n 0.0113869f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_200 VPB N_D_M1005_g 0.0397993f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.16
cc_201 VPB D 0.00128041f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.805
cc_202 VPB N_D_c_392_n 0.0257434f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.885
cc_203 VPB N_A_332_93#_M1041_g 0.0248503f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.16
cc_204 VPB N_A_332_93#_c_442_n 0.0187025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_332_93#_c_443_n 0.0241887f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_206 VPB N_A_332_93#_c_437_n 0.00520453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_332_93#_c_445_n 0.00828601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_332_93#_c_446_n 0.0148647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_332_93#_c_439_n 0.0119623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_332_93#_c_440_n 0.027809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_332_93#_c_449_n 0.00548065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_SCE_M1032_g 0.0204979f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.805
cc_213 VPB N_SCE_M1038_g 0.0292204f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_214 VPB N_SCE_c_535_n 0.0119814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_SCE_c_536_n 0.00930402f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.55
cc_216 VPB N_SCE_c_530_n 0.0286079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_SCE_c_538_n 0.0131628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB SCE 0.00481753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_SCE_c_532_n 0.017024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_CLK_M1006_g 0.0292326f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.16
cc_221 VPB N_CLK_c_625_n 0.0293585f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.16
cc_222 VPB N_CLK_c_626_n 0.0378783f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.72
cc_223 VPB CLK 0.00624387f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.12
cc_224 VPB N_CLK_c_623_n 7.68063e-19 $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_225 VPB N_A_893_101#_M1012_g 0.0500236f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.31
cc_226 VPB N_A_893_101#_c_681_n 0.0615229f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_227 VPB N_A_893_101#_c_672_n 0.00533665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_893_101#_c_683_n 0.0110478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_893_101#_c_684_n 0.00246661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_893_101#_c_685_n 0.00825021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_893_101#_c_686_n 0.00536992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_893_101#_c_676_n 0.0366198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_893_101#_c_677_n 0.0152025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_893_101#_c_679_n 0.00369993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_1297_290#_M1016_g 0.0422619f $X=-0.19 $Y=1.655 $X2=0.555
+ $Y2=0.805
cc_236 VPB N_A_1297_290#_M1031_g 0.0207038f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.27
cc_237 VPB N_A_1297_290#_c_839_n 0.00518703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_1297_290#_c_840_n 7.12703e-19 $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.38
cc_239 VPB N_A_1297_290#_c_851_n 0.00610718f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.55
cc_240 VPB N_A_1297_290#_c_852_n 0.00240335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_1297_290#_c_842_n 0.00198494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1297_290#_c_854_n 0.00421873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1297_290#_c_843_n 0.0039035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1297_290#_c_844_n 0.00472013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_1297_290#_c_845_n 7.98646e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1297_290#_c_846_n 0.0180665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_SET_B_M1040_g 0.0188243f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.16
cc_248 VPB N_SET_B_M1011_g 0.00374028f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.31
cc_249 VPB N_SET_B_c_1019_n 0.0252695f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.31
cc_250 VPB N_SET_B_M1020_g 0.0225239f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.885
cc_251 VPB N_SET_B_c_1027_n 0.00189137f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_252 VPB SET_B 0.00459914f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_SET_B_c_1029_n 0.0152707f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_254 VPB N_SET_B_c_1030_n 0.00133112f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_255 VPB N_SET_B_c_1021_n 0.00130945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_SET_B_c_1022_n 0.00806029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_SET_B_c_1033_n 0.00324263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_SET_B_c_1034_n 0.00123149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_1216_457#_M1024_g 0.0192968f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.31
cc_260 VPB N_A_1216_457#_c_1155_n 0.00784301f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_261 VPB N_A_1216_457#_c_1157_n 0.0136757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_1216_457#_c_1160_n 0.00127954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_1650_21#_M1046_g 0.0194575f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.16
cc_264 VPB N_A_1650_21#_M1014_g 0.0247451f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.12
cc_265 VPB N_A_1650_21#_c_1252_n 0.0206173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_1650_21#_c_1263_n 0.0183823f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_755_106#_M1042_g 0.0510843f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.885
cc_268 VPB N_A_755_106#_c_1436_n 0.102896f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_269 VPB N_A_755_106#_c_1437_n 0.012806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_755_106#_M1043_g 0.0417059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_755_106#_c_1439_n 0.211474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_755_106#_M1035_g 0.00992761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_755_106#_c_1441_n 0.0478121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_755_106#_c_1442_n 0.0416247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_755_106#_M1027_g 0.00197417f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_755_106#_c_1444_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_755_106#_c_1433_n 0.0147155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_755_106#_c_1446_n 0.0240452f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_755_106#_c_1434_n 0.00314273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_2064_453#_M1017_g 0.0251187f $X=-0.19 $Y=1.655 $X2=0.555
+ $Y2=0.805
cc_281 VPB N_A_2064_453#_M1009_g 0.00538603f $X=-0.19 $Y=1.655 $X2=0.425
+ $Y2=1.31
cc_282 VPB N_A_2064_453#_M1045_g 0.0254051f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_283 VPB N_A_2064_453#_M1025_g 0.0257557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_2064_453#_c_1596_n 0.0633357f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_A_2064_453#_c_1597_n 0.00154871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_A_2064_453#_c_1598_n 0.0169139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_A_2064_453#_c_1599_n 0.0044134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_A_2064_453#_c_1600_n 0.00648746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_A_2064_453#_c_1587_n 0.0017335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_A_2064_453#_c_1602_n 0.0157427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_A_2064_453#_c_1588_n 0.0017426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_A_1861_431#_M1021_g 0.021266f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.31
cc_293 VPB N_A_1861_431#_c_1756_n 0.00948356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_A_1861_431#_c_1764_n 0.00271415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_RESET_B_M1000_g 0.0258832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_A_2892_137#_M1044_g 0.0281256f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.31
cc_297 VPB N_A_2892_137#_c_1915_n 0.00649261f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.38
cc_298 VPB N_A_27_481#_c_1960_n 0.0343396f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.805
cc_299 VPB N_A_27_481#_c_1961_n 0.0173163f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.31
cc_300 VPB N_A_27_481#_c_1962_n 0.0100305f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.16
cc_301 VPB N_A_27_481#_c_1963_n 0.0025298f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.72
cc_302 VPB N_A_27_481#_c_1964_n 0.00690381f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.885
cc_303 VPB N_A_27_481#_c_1965_n 0.00140515f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.12
cc_304 VPB N_A_27_481#_c_1966_n 0.00852962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_2011_n 0.00711854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2012_n 0.0163577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2013_n 0.0204586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2014_n 0.0134734f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2015_n 0.0222444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2016_n 0.0153388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2017_n 0.0122469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2018_n 0.00434291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2019_n 0.018542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_2020_n 0.0193798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_2021_n 0.0176719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_2022_n 0.0306876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_2023_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_2024_n 0.0275934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_2025_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_2026_n 0.0331938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_2027_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_2028_n 0.019006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_2029_n 0.0398854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_2030_n 0.0457779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2031_n 0.0309695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_2032_n 0.0654578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_2033_n 0.0238029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2034_n 0.0191143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_2010_n 0.14743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_2036_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2037_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_2038_n 0.00575291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_2039_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2040_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_2041_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_2042_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_A_204_119#_c_2218_n 5.94466e-19 $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.38
cc_338 VPB N_A_204_119#_c_2202_n 0.00349683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_A_204_119#_c_2220_n 0.0088519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_A_204_119#_c_2221_n 0.0103478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_A_204_119#_c_2216_n 0.0090451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_342 VPB N_Q_N_c_2398_n 0.00481231f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.12
cc_343 VPB N_Q_N_c_2397_n 0.00305494f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.27
cc_344 VPB Q_N 0.0210645f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_345 VPB N_Q_c_2432_n 0.0429721f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.805
cc_346 VPB N_Q_c_2433_n 0.0137223f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.72
cc_347 VPB N_Q_c_2429_n 0.00779836f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.885
cc_348 N_SCD_M1033_g N_SCE_M1013_g 0.0429225f $X=0.555 $Y=0.805 $X2=0 $Y2=0
cc_349 N_SCD_c_351_n N_SCE_M1013_g 0.00841712f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_350 N_SCD_c_352_n N_SCE_M1013_g 0.00165586f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_351 N_SCD_c_356_n N_SCE_M1032_g 0.0172793f $X=0.485 $Y=2.27 $X2=0 $Y2=0
cc_352 N_SCD_c_354_n N_SCE_c_535_n 0.00423555f $X=0.385 $Y=1.885 $X2=0 $Y2=0
cc_353 N_SCD_c_355_n N_SCE_c_536_n 0.00423555f $X=0.485 $Y=2.12 $X2=0 $Y2=0
cc_354 N_SCD_c_356_n N_SCE_c_536_n 0.00388451f $X=0.485 $Y=2.27 $X2=0 $Y2=0
cc_355 N_SCD_c_351_n SCE 4.11905e-19 $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_356 N_SCD_c_352_n SCE 0.0221109f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_357 N_SCD_c_351_n N_SCE_c_532_n 0.0213895f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_358 N_SCD_c_352_n N_SCE_c_532_n 4.12997e-19 $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_359 N_SCD_M1037_g N_A_27_481#_c_1960_n 0.0130012f $X=0.495 $Y=2.725 $X2=0
+ $Y2=0
cc_360 N_SCD_c_356_n N_A_27_481#_c_1960_n 0.00192345f $X=0.485 $Y=2.27 $X2=0
+ $Y2=0
cc_361 N_SCD_c_355_n N_A_27_481#_c_1961_n 0.00278222f $X=0.485 $Y=2.12 $X2=0
+ $Y2=0
cc_362 N_SCD_c_356_n N_A_27_481#_c_1961_n 0.00877399f $X=0.485 $Y=2.27 $X2=0
+ $Y2=0
cc_363 N_SCD_c_352_n N_A_27_481#_c_1961_n 0.00756021f $X=0.385 $Y=1.38 $X2=0
+ $Y2=0
cc_364 N_SCD_c_354_n N_A_27_481#_c_1962_n 0.00487488f $X=0.385 $Y=1.885 $X2=0
+ $Y2=0
cc_365 N_SCD_c_355_n N_A_27_481#_c_1962_n 0.00197483f $X=0.485 $Y=2.12 $X2=0
+ $Y2=0
cc_366 N_SCD_c_356_n N_A_27_481#_c_1962_n 0.00277464f $X=0.485 $Y=2.27 $X2=0
+ $Y2=0
cc_367 N_SCD_c_352_n N_A_27_481#_c_1962_n 0.0273972f $X=0.385 $Y=1.38 $X2=0
+ $Y2=0
cc_368 N_SCD_M1037_g N_VPWR_c_2011_n 0.00642796f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_369 N_SCD_M1037_g N_VPWR_c_2028_n 0.00502664f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_370 N_SCD_M1037_g N_VPWR_c_2010_n 0.0102756f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_371 N_SCD_M1033_g N_A_204_119#_c_2199_n 0.00199884f $X=0.555 $Y=0.805 $X2=0
+ $Y2=0
cc_372 N_SCD_c_350_n N_A_204_119#_c_2201_n 5.30423e-19 $X=0.425 $Y=1.31 $X2=0
+ $Y2=0
cc_373 N_SCD_c_352_n N_A_204_119#_c_2201_n 0.00479053f $X=0.385 $Y=1.38 $X2=0
+ $Y2=0
cc_374 N_SCD_M1033_g N_VGND_c_2455_n 0.0141328f $X=0.555 $Y=0.805 $X2=0 $Y2=0
cc_375 N_SCD_c_350_n N_VGND_c_2455_n 0.00751937f $X=0.425 $Y=1.31 $X2=0 $Y2=0
cc_376 N_SCD_c_352_n N_VGND_c_2455_n 0.0279363f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_377 N_SCD_M1033_g N_VGND_c_2464_n 0.0035863f $X=0.555 $Y=0.805 $X2=0 $Y2=0
cc_378 N_SCD_M1033_g N_VGND_c_2480_n 0.00401353f $X=0.555 $Y=0.805 $X2=0 $Y2=0
cc_379 N_D_M1019_g N_A_332_93#_c_433_n 0.0462106f $X=1.375 $Y=0.805 $X2=0 $Y2=0
cc_380 N_D_c_392_n N_A_332_93#_c_435_n 0.0055001f $X=1.625 $Y=1.69 $X2=0 $Y2=0
cc_381 N_D_M1019_g N_A_332_93#_c_436_n 0.00317896f $X=1.375 $Y=0.805 $X2=0 $Y2=0
cc_382 N_D_M1005_g N_A_332_93#_c_442_n 0.0028982f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_383 N_D_M1005_g N_A_332_93#_c_443_n 0.0334694f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_384 D N_A_332_93#_c_437_n 0.00103106f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_385 N_D_c_392_n N_A_332_93#_c_437_n 0.0215456f $X=1.625 $Y=1.69 $X2=0 $Y2=0
cc_386 N_D_M1019_g N_SCE_M1013_g 0.0330782f $X=1.375 $Y=0.805 $X2=0 $Y2=0
cc_387 N_D_M1019_g N_SCE_c_525_n 0.0103003f $X=1.375 $Y=0.805 $X2=0 $Y2=0
cc_388 N_D_M1005_g N_SCE_c_536_n 0.0501906f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_389 N_D_M1005_g SCE 6.89287e-19 $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_390 D SCE 0.0240649f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_391 N_D_c_392_n SCE 0.00268301f $X=1.625 $Y=1.69 $X2=0 $Y2=0
cc_392 N_D_M1005_g N_SCE_c_532_n 0.0118204f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_393 D N_SCE_c_532_n 2.10045e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_394 N_D_c_392_n N_SCE_c_532_n 0.0193616f $X=1.625 $Y=1.69 $X2=0 $Y2=0
cc_395 N_D_M1005_g N_A_27_481#_c_1961_n 0.00134936f $X=1.435 $Y=2.725 $X2=0
+ $Y2=0
cc_396 N_D_c_392_n N_A_27_481#_c_1961_n 2.31726e-19 $X=1.625 $Y=1.69 $X2=0 $Y2=0
cc_397 N_D_M1005_g N_A_27_481#_c_1963_n 0.00291362f $X=1.435 $Y=2.725 $X2=0
+ $Y2=0
cc_398 N_D_M1005_g N_A_27_481#_c_1964_n 0.0127852f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_399 N_D_M1005_g N_VPWR_c_2029_n 0.00327726f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_400 N_D_M1005_g N_VPWR_c_2010_n 0.004836f $X=1.435 $Y=2.725 $X2=0 $Y2=0
cc_401 N_D_M1019_g N_A_204_119#_c_2199_n 0.0125542f $X=1.375 $Y=0.805 $X2=0
+ $Y2=0
cc_402 N_D_M1019_g N_A_204_119#_c_2200_n 0.0158499f $X=1.375 $Y=0.805 $X2=0
+ $Y2=0
cc_403 D N_A_204_119#_c_2200_n 0.023777f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_404 N_D_c_392_n N_A_204_119#_c_2200_n 0.00594777f $X=1.625 $Y=1.69 $X2=0
+ $Y2=0
cc_405 N_D_M1019_g N_A_204_119#_c_2201_n 0.00360577f $X=1.375 $Y=0.805 $X2=0
+ $Y2=0
cc_406 N_D_M1005_g N_A_204_119#_c_2218_n 0.00797403f $X=1.435 $Y=2.725 $X2=0
+ $Y2=0
cc_407 N_D_M1019_g N_A_204_119#_c_2202_n 0.00272615f $X=1.375 $Y=0.805 $X2=0
+ $Y2=0
cc_408 N_D_M1005_g N_A_204_119#_c_2202_n 0.0031372f $X=1.435 $Y=2.725 $X2=0
+ $Y2=0
cc_409 D N_A_204_119#_c_2202_n 0.0250785f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_410 N_D_c_392_n N_A_204_119#_c_2202_n 9.58437e-19 $X=1.625 $Y=1.69 $X2=0
+ $Y2=0
cc_411 N_D_M1005_g N_A_204_119#_c_2220_n 0.00512686f $X=1.435 $Y=2.725 $X2=0
+ $Y2=0
cc_412 D N_A_204_119#_c_2220_n 0.0222428f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_413 N_D_c_392_n N_A_204_119#_c_2220_n 0.00623744f $X=1.625 $Y=1.69 $X2=0
+ $Y2=0
cc_414 N_D_M1019_g N_VGND_c_2456_n 0.0016998f $X=1.375 $Y=0.805 $X2=0 $Y2=0
cc_415 N_D_M1019_g N_VGND_c_2480_n 9.39239e-19 $X=1.375 $Y=0.805 $X2=0 $Y2=0
cc_416 N_A_332_93#_c_433_n N_SCE_c_525_n 0.0103107f $X=1.735 $Y=1.09 $X2=0 $Y2=0
cc_417 N_A_332_93#_c_433_n N_SCE_M1034_g 0.0069113f $X=1.735 $Y=1.09 $X2=0 $Y2=0
cc_418 N_A_332_93#_c_438_n N_SCE_M1034_g 0.00192143f $X=2.65 $Y=0.825 $X2=0
+ $Y2=0
cc_419 N_A_332_93#_c_438_n N_SCE_c_528_n 0.0130924f $X=2.65 $Y=0.825 $X2=0 $Y2=0
cc_420 N_A_332_93#_c_445_n N_SCE_c_528_n 0.00408667f $X=2.985 $Y=1.77 $X2=0
+ $Y2=0
cc_421 N_A_332_93#_c_434_n N_SCE_c_529_n 0.0096783f $X=2 $Y=1.165 $X2=0 $Y2=0
cc_422 N_A_332_93#_c_439_n N_SCE_c_529_n 0.00129657f $X=2.49 $Y=1.69 $X2=0 $Y2=0
cc_423 N_A_332_93#_c_440_n N_SCE_c_529_n 0.0130384f $X=2.49 $Y=1.69 $X2=0 $Y2=0
cc_424 N_A_332_93#_c_446_n N_SCE_M1038_g 0.00836774f $X=3.15 $Y=2.55 $X2=0 $Y2=0
cc_425 N_A_332_93#_c_449_n N_SCE_M1038_g 0.00794832f $X=3.15 $Y=2.385 $X2=0
+ $Y2=0
cc_426 N_A_332_93#_c_438_n N_SCE_c_530_n 0.0125469f $X=2.65 $Y=0.825 $X2=0 $Y2=0
cc_427 N_A_332_93#_c_445_n N_SCE_c_530_n 0.0125187f $X=2.985 $Y=1.77 $X2=0 $Y2=0
cc_428 N_A_332_93#_c_440_n N_SCE_c_530_n 0.0173388f $X=2.49 $Y=1.69 $X2=0 $Y2=0
cc_429 N_A_332_93#_c_449_n N_SCE_c_530_n 0.0123887f $X=3.15 $Y=2.385 $X2=0 $Y2=0
cc_430 N_A_332_93#_c_443_n N_SCE_c_538_n 0.00348722f $X=2.075 $Y=2.17 $X2=0
+ $Y2=0
cc_431 N_A_332_93#_c_445_n N_SCE_c_538_n 0.0013475f $X=2.985 $Y=1.77 $X2=0 $Y2=0
cc_432 N_A_332_93#_c_449_n N_SCE_c_538_n 0.00932532f $X=3.15 $Y=2.385 $X2=0
+ $Y2=0
cc_433 N_A_332_93#_c_446_n N_CLK_M1006_g 0.00129898f $X=3.15 $Y=2.55 $X2=0 $Y2=0
cc_434 N_A_332_93#_c_449_n N_CLK_M1006_g 0.00368033f $X=3.15 $Y=2.385 $X2=0
+ $Y2=0
cc_435 N_A_332_93#_c_445_n N_CLK_c_625_n 0.00133744f $X=2.985 $Y=1.77 $X2=0
+ $Y2=0
cc_436 N_A_332_93#_c_449_n N_CLK_c_625_n 0.00234313f $X=3.15 $Y=2.385 $X2=0
+ $Y2=0
cc_437 N_A_332_93#_c_445_n CLK 0.00925756f $X=2.985 $Y=1.77 $X2=0 $Y2=0
cc_438 N_A_332_93#_c_449_n CLK 0.0158428f $X=3.15 $Y=2.385 $X2=0 $Y2=0
cc_439 N_A_332_93#_M1041_g N_A_27_481#_c_1964_n 0.0150064f $X=1.865 $Y=2.725
+ $X2=0 $Y2=0
cc_440 N_A_332_93#_M1041_g N_A_27_481#_c_1966_n 0.00983386f $X=1.865 $Y=2.725
+ $X2=0 $Y2=0
cc_441 N_A_332_93#_c_443_n N_A_27_481#_c_1966_n 0.00444387f $X=2.075 $Y=2.17
+ $X2=0 $Y2=0
cc_442 N_A_332_93#_c_440_n N_A_27_481#_c_1966_n 0.00525575f $X=2.49 $Y=1.69
+ $X2=0 $Y2=0
cc_443 N_A_332_93#_M1041_g N_VPWR_c_2012_n 0.00290616f $X=1.865 $Y=2.725 $X2=0
+ $Y2=0
cc_444 N_A_332_93#_c_445_n N_VPWR_c_2012_n 0.00264375f $X=2.985 $Y=1.77 $X2=0
+ $Y2=0
cc_445 N_A_332_93#_c_446_n N_VPWR_c_2012_n 0.0257922f $X=3.15 $Y=2.55 $X2=0
+ $Y2=0
cc_446 N_A_332_93#_c_439_n N_VPWR_c_2012_n 0.00707052f $X=2.49 $Y=1.69 $X2=0
+ $Y2=0
cc_447 N_A_332_93#_c_440_n N_VPWR_c_2012_n 6.51034e-19 $X=2.49 $Y=1.69 $X2=0
+ $Y2=0
cc_448 N_A_332_93#_c_446_n N_VPWR_c_2013_n 0.0220321f $X=3.15 $Y=2.55 $X2=0
+ $Y2=0
cc_449 N_A_332_93#_c_446_n N_VPWR_c_2014_n 0.0458108f $X=3.15 $Y=2.55 $X2=0
+ $Y2=0
cc_450 N_A_332_93#_c_449_n N_VPWR_c_2014_n 0.00154216f $X=3.15 $Y=2.385 $X2=0
+ $Y2=0
cc_451 N_A_332_93#_M1041_g N_VPWR_c_2029_n 0.00327726f $X=1.865 $Y=2.725 $X2=0
+ $Y2=0
cc_452 N_A_332_93#_M1041_g N_VPWR_c_2010_n 0.00578801f $X=1.865 $Y=2.725 $X2=0
+ $Y2=0
cc_453 N_A_332_93#_c_446_n N_VPWR_c_2010_n 0.0125808f $X=3.15 $Y=2.55 $X2=0
+ $Y2=0
cc_454 N_A_332_93#_c_433_n N_A_204_119#_c_2199_n 0.00209048f $X=1.735 $Y=1.09
+ $X2=0 $Y2=0
cc_455 N_A_332_93#_c_434_n N_A_204_119#_c_2200_n 0.00489152f $X=2 $Y=1.165 $X2=0
+ $Y2=0
cc_456 N_A_332_93#_c_435_n N_A_204_119#_c_2200_n 0.00854778f $X=1.81 $Y=1.165
+ $X2=0 $Y2=0
cc_457 N_A_332_93#_M1041_g N_A_204_119#_c_2218_n 0.0118177f $X=1.865 $Y=2.725
+ $X2=0 $Y2=0
cc_458 N_A_332_93#_c_443_n N_A_204_119#_c_2218_n 0.00238135f $X=2.075 $Y=2.17
+ $X2=0 $Y2=0
cc_459 N_A_332_93#_c_436_n N_A_204_119#_c_2202_n 0.00689279f $X=2.075 $Y=1.525
+ $X2=0 $Y2=0
cc_460 N_A_332_93#_c_442_n N_A_204_119#_c_2202_n 0.0109997f $X=2.075 $Y=2.095
+ $X2=0 $Y2=0
cc_461 N_A_332_93#_c_443_n N_A_204_119#_c_2202_n 2.07993e-19 $X=2.075 $Y=2.17
+ $X2=0 $Y2=0
cc_462 N_A_332_93#_c_437_n N_A_204_119#_c_2202_n 0.00974802f $X=2.075 $Y=1.69
+ $X2=0 $Y2=0
cc_463 N_A_332_93#_c_438_n N_A_204_119#_c_2202_n 0.00652736f $X=2.65 $Y=0.825
+ $X2=0 $Y2=0
cc_464 N_A_332_93#_c_439_n N_A_204_119#_c_2202_n 0.0229098f $X=2.49 $Y=1.69
+ $X2=0 $Y2=0
cc_465 N_A_332_93#_c_433_n N_A_204_119#_c_2203_n 0.00255854f $X=1.735 $Y=1.09
+ $X2=0 $Y2=0
cc_466 N_A_332_93#_c_434_n N_A_204_119#_c_2203_n 0.00200718f $X=2 $Y=1.165 $X2=0
+ $Y2=0
cc_467 N_A_332_93#_c_438_n N_A_204_119#_c_2203_n 0.0235215f $X=2.65 $Y=0.825
+ $X2=0 $Y2=0
cc_468 N_A_332_93#_c_438_n N_A_204_119#_c_2204_n 0.0123913f $X=2.65 $Y=0.825
+ $X2=0 $Y2=0
cc_469 N_A_332_93#_c_438_n N_A_204_119#_c_2206_n 0.0376637f $X=2.65 $Y=0.825
+ $X2=0 $Y2=0
cc_470 N_A_332_93#_c_445_n N_A_204_119#_c_2207_n 0.00345632f $X=2.985 $Y=1.77
+ $X2=0 $Y2=0
cc_471 N_A_332_93#_c_438_n N_A_204_119#_c_2208_n 0.0126276f $X=2.65 $Y=0.825
+ $X2=0 $Y2=0
cc_472 N_A_332_93#_c_445_n N_A_204_119#_c_2208_n 0.00779738f $X=2.985 $Y=1.77
+ $X2=0 $Y2=0
cc_473 N_A_332_93#_c_442_n N_A_204_119#_c_2220_n 0.00373222f $X=2.075 $Y=2.095
+ $X2=0 $Y2=0
cc_474 N_A_332_93#_c_443_n N_A_204_119#_c_2220_n 0.0214693f $X=2.075 $Y=2.17
+ $X2=0 $Y2=0
cc_475 N_A_332_93#_c_434_n N_A_204_119#_c_2215_n 0.00681281f $X=2 $Y=1.165 $X2=0
+ $Y2=0
cc_476 N_A_332_93#_c_436_n N_A_204_119#_c_2215_n 0.00439412f $X=2.075 $Y=1.525
+ $X2=0 $Y2=0
cc_477 N_A_332_93#_c_438_n N_A_204_119#_c_2215_n 0.0130902f $X=2.65 $Y=0.825
+ $X2=0 $Y2=0
cc_478 N_A_332_93#_c_439_n N_A_204_119#_c_2215_n 0.00426713f $X=2.49 $Y=1.69
+ $X2=0 $Y2=0
cc_479 N_A_332_93#_c_440_n N_A_204_119#_c_2215_n 0.00683719f $X=2.49 $Y=1.69
+ $X2=0 $Y2=0
cc_480 N_A_332_93#_c_433_n N_VGND_c_2456_n 0.0111257f $X=1.735 $Y=1.09 $X2=0
+ $Y2=0
cc_481 N_A_332_93#_c_434_n N_VGND_c_2456_n 0.00496753f $X=2 $Y=1.165 $X2=0 $Y2=0
cc_482 N_A_332_93#_c_433_n N_VGND_c_2480_n 7.88961e-19 $X=1.735 $Y=1.09 $X2=0
+ $Y2=0
cc_483 N_SCE_c_528_n N_CLK_M1015_g 0.00802767f $X=2.895 $Y=1.165 $X2=0 $Y2=0
cc_484 N_SCE_c_538_n N_CLK_c_625_n 0.00959488f $X=2.952 $Y=2.245 $X2=0 $Y2=0
cc_485 N_SCE_c_530_n CLK 0.00159511f $X=2.952 $Y=2.095 $X2=0 $Y2=0
cc_486 N_SCE_c_530_n N_CLK_c_623_n 0.00959488f $X=2.952 $Y=2.095 $X2=0 $Y2=0
cc_487 N_SCE_M1032_g N_A_27_481#_c_1960_n 9.22263e-19 $X=1.045 $Y=2.725 $X2=0
+ $Y2=0
cc_488 N_SCE_c_535_n N_A_27_481#_c_1961_n 0.00320334f $X=1.03 $Y=2.095 $X2=0
+ $Y2=0
cc_489 N_SCE_c_536_n N_A_27_481#_c_1961_n 0.0131211f $X=1.03 $Y=2.245 $X2=0
+ $Y2=0
cc_490 SCE N_A_27_481#_c_1961_n 0.0385273f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_491 N_SCE_c_532_n N_A_27_481#_c_1961_n 0.00426808f $X=0.925 $Y=1.715 $X2=0
+ $Y2=0
cc_492 N_SCE_c_536_n N_A_27_481#_c_1963_n 0.00608438f $X=1.03 $Y=2.245 $X2=0
+ $Y2=0
cc_493 N_SCE_M1032_g N_A_27_481#_c_1965_n 7.64437e-19 $X=1.045 $Y=2.725 $X2=0
+ $Y2=0
cc_494 N_SCE_M1032_g N_VPWR_c_2011_n 0.00453029f $X=1.045 $Y=2.725 $X2=0 $Y2=0
cc_495 N_SCE_M1038_g N_VPWR_c_2012_n 0.00476117f $X=2.935 $Y=2.725 $X2=0 $Y2=0
cc_496 N_SCE_M1038_g N_VPWR_c_2013_n 0.00502664f $X=2.935 $Y=2.725 $X2=0 $Y2=0
cc_497 N_SCE_M1038_g N_VPWR_c_2014_n 0.00329606f $X=2.935 $Y=2.725 $X2=0 $Y2=0
cc_498 N_SCE_M1032_g N_VPWR_c_2029_n 0.0053602f $X=1.045 $Y=2.725 $X2=0 $Y2=0
cc_499 N_SCE_M1032_g N_VPWR_c_2010_n 0.0103449f $X=1.045 $Y=2.725 $X2=0 $Y2=0
cc_500 N_SCE_M1038_g N_VPWR_c_2010_n 0.011218f $X=2.935 $Y=2.725 $X2=0 $Y2=0
cc_501 N_SCE_M1013_g N_A_204_119#_c_2199_n 0.0130485f $X=0.945 $Y=0.805 $X2=0
+ $Y2=0
cc_502 N_SCE_c_525_n N_A_204_119#_c_2199_n 0.00392786f $X=2.36 $Y=0.18 $X2=0
+ $Y2=0
cc_503 N_SCE_M1013_g N_A_204_119#_c_2201_n 0.0052373f $X=0.945 $Y=0.805 $X2=0
+ $Y2=0
cc_504 SCE N_A_204_119#_c_2201_n 0.0219628f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_505 N_SCE_c_532_n N_A_204_119#_c_2201_n 0.00186749f $X=0.925 $Y=1.715 $X2=0
+ $Y2=0
cc_506 N_SCE_M1034_g N_A_204_119#_c_2203_n 0.0167848f $X=2.435 $Y=0.805 $X2=0
+ $Y2=0
cc_507 N_SCE_c_529_n N_A_204_119#_c_2203_n 0.00193042f $X=2.51 $Y=1.165 $X2=0
+ $Y2=0
cc_508 N_SCE_M1034_g N_A_204_119#_c_2204_n 0.0124521f $X=2.435 $Y=0.805 $X2=0
+ $Y2=0
cc_509 N_SCE_c_528_n N_A_204_119#_c_2204_n 0.00544133f $X=2.895 $Y=1.165 $X2=0
+ $Y2=0
cc_510 N_SCE_c_525_n N_A_204_119#_c_2205_n 0.00135484f $X=2.36 $Y=0.18 $X2=0
+ $Y2=0
cc_511 N_SCE_M1034_g N_A_204_119#_c_2205_n 0.00355912f $X=2.435 $Y=0.805 $X2=0
+ $Y2=0
cc_512 N_SCE_M1034_g N_A_204_119#_c_2206_n 0.00377575f $X=2.435 $Y=0.805 $X2=0
+ $Y2=0
cc_513 N_SCE_c_528_n N_A_204_119#_c_2206_n 0.00535238f $X=2.895 $Y=1.165 $X2=0
+ $Y2=0
cc_514 N_SCE_c_528_n N_A_204_119#_c_2208_n 0.00418411f $X=2.895 $Y=1.165 $X2=0
+ $Y2=0
cc_515 N_SCE_c_530_n N_A_204_119#_c_2208_n 0.00578315f $X=2.952 $Y=2.095 $X2=0
+ $Y2=0
cc_516 N_SCE_c_528_n N_A_204_119#_c_2209_n 2.1243e-19 $X=2.895 $Y=1.165 $X2=0
+ $Y2=0
cc_517 N_SCE_c_529_n N_A_204_119#_c_2215_n 0.00192721f $X=2.51 $Y=1.165 $X2=0
+ $Y2=0
cc_518 N_SCE_M1013_g N_VGND_c_2455_n 0.0018473f $X=0.945 $Y=0.805 $X2=0 $Y2=0
cc_519 N_SCE_c_526_n N_VGND_c_2455_n 0.00977077f $X=1.02 $Y=0.18 $X2=0 $Y2=0
cc_520 N_SCE_c_525_n N_VGND_c_2456_n 0.0210723f $X=2.36 $Y=0.18 $X2=0 $Y2=0
cc_521 N_SCE_M1034_g N_VGND_c_2456_n 0.00286637f $X=2.435 $Y=0.805 $X2=0 $Y2=0
cc_522 N_SCE_c_526_n N_VGND_c_2464_n 0.0294461f $X=1.02 $Y=0.18 $X2=0 $Y2=0
cc_523 N_SCE_c_525_n N_VGND_c_2466_n 0.0131867f $X=2.36 $Y=0.18 $X2=0 $Y2=0
cc_524 N_SCE_c_525_n N_VGND_c_2480_n 0.0465559f $X=2.36 $Y=0.18 $X2=0 $Y2=0
cc_525 N_SCE_c_526_n N_VGND_c_2480_n 0.0107881f $X=1.02 $Y=0.18 $X2=0 $Y2=0
cc_526 N_CLK_M1015_g N_A_755_106#_c_1422_n 0.0186386f $X=3.7 $Y=0.74 $X2=0 $Y2=0
cc_527 N_CLK_M1015_g N_A_755_106#_c_1432_n 0.00681535f $X=3.7 $Y=0.74 $X2=0
+ $Y2=0
cc_528 CLK N_A_755_106#_c_1432_n 0.0168627f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_529 CLK N_A_755_106#_c_1433_n 2.68148e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_530 N_CLK_c_623_n N_A_755_106#_c_1433_n 0.0186386f $X=3.61 $Y=1.665 $X2=0
+ $Y2=0
cc_531 N_CLK_c_625_n N_A_755_106#_c_1446_n 0.00611045f $X=3.61 $Y=2.02 $X2=0
+ $Y2=0
cc_532 N_CLK_c_626_n N_A_755_106#_c_1446_n 0.0129316f $X=3.925 $Y=2.095 $X2=0
+ $Y2=0
cc_533 CLK N_A_755_106#_c_1446_n 0.0237138f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_534 N_CLK_c_626_n N_A_755_106#_c_1434_n 0.00144695f $X=3.925 $Y=2.095 $X2=0
+ $Y2=0
cc_535 N_CLK_c_623_n N_A_755_106#_c_1434_n 0.00279263f $X=3.61 $Y=1.665 $X2=0
+ $Y2=0
cc_536 N_CLK_M1006_g N_VPWR_c_2014_n 0.015593f $X=3.925 $Y=2.69 $X2=0 $Y2=0
cc_537 N_CLK_c_626_n N_VPWR_c_2014_n 0.00486883f $X=3.925 $Y=2.095 $X2=0 $Y2=0
cc_538 CLK N_VPWR_c_2014_n 0.019442f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_539 N_CLK_M1006_g N_VPWR_c_2022_n 0.00418439f $X=3.925 $Y=2.69 $X2=0 $Y2=0
cc_540 N_CLK_M1006_g N_VPWR_c_2010_n 0.00845728f $X=3.925 $Y=2.69 $X2=0 $Y2=0
cc_541 N_CLK_M1015_g N_A_204_119#_c_2206_n 0.00148593f $X=3.7 $Y=0.74 $X2=0
+ $Y2=0
cc_542 N_CLK_M1015_g N_A_204_119#_c_2207_n 0.00822553f $X=3.7 $Y=0.74 $X2=0
+ $Y2=0
cc_543 N_CLK_c_626_n N_A_204_119#_c_2207_n 2.38481e-19 $X=3.925 $Y=2.095 $X2=0
+ $Y2=0
cc_544 CLK N_A_204_119#_c_2207_n 0.0257599f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_545 N_CLK_c_623_n N_A_204_119#_c_2207_n 0.00123812f $X=3.61 $Y=1.665 $X2=0
+ $Y2=0
cc_546 N_CLK_M1015_g N_A_204_119#_c_2209_n 0.0281954f $X=3.7 $Y=0.74 $X2=0 $Y2=0
cc_547 N_CLK_M1015_g N_A_204_119#_c_2211_n 0.00438273f $X=3.7 $Y=0.74 $X2=0
+ $Y2=0
cc_548 N_CLK_M1015_g N_VGND_c_2457_n 0.00392799f $X=3.7 $Y=0.74 $X2=0 $Y2=0
cc_549 N_CLK_M1015_g N_VGND_c_2468_n 6.68053e-19 $X=3.7 $Y=0.74 $X2=0 $Y2=0
cc_550 N_A_893_101#_M1012_g N_A_1297_290#_M1016_g 0.00328955f $X=6.005 $Y=2.495
+ $X2=0 $Y2=0
cc_551 N_A_893_101#_c_665_n N_A_1297_290#_M1010_g 0.00256418f $X=6.005 $Y=1.415
+ $X2=0 $Y2=0
cc_552 N_A_893_101#_c_667_n N_A_1297_290#_M1010_g 0.00155541f $X=6.37 $Y=1.165
+ $X2=0 $Y2=0
cc_553 N_A_893_101#_M1023_g N_A_1297_290#_M1010_g 0.0673073f $X=6.515 $Y=0.445
+ $X2=0 $Y2=0
cc_554 N_A_893_101#_c_673_n N_A_1297_290#_M1010_g 0.00660819f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_555 N_A_893_101#_c_673_n N_A_1297_290#_c_840_n 0.00637292f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_556 N_A_893_101#_M1018_g N_A_1297_290#_M1008_g 0.0418279f $X=9.745 $Y=0.605
+ $X2=0 $Y2=0
cc_557 N_A_893_101#_c_673_n N_A_1297_290#_c_866_n 0.006879f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_558 N_A_893_101#_c_673_n N_A_1297_290#_c_867_n 0.00612926f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_559 N_A_893_101#_c_673_n N_A_1297_290#_c_842_n 0.0179675f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_560 N_A_893_101#_c_673_n N_A_1297_290#_c_854_n 0.0171033f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_561 N_A_893_101#_c_679_n N_A_1297_290#_c_854_n 0.00864363f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_562 N_A_893_101#_c_673_n N_A_1297_290#_c_843_n 0.0259679f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_563 N_A_893_101#_c_675_n N_A_1297_290#_c_843_n 5.25698e-19 $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_564 N_A_893_101#_c_678_n N_A_1297_290#_c_843_n 0.00107576f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_565 N_A_893_101#_c_679_n N_A_1297_290#_c_843_n 0.0472168f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_566 N_A_893_101#_c_673_n N_A_1297_290#_c_844_n 0.00282036f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_567 N_A_893_101#_c_678_n N_A_1297_290#_c_844_n 0.0217086f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_568 N_A_893_101#_c_679_n N_A_1297_290#_c_844_n 0.00227336f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_569 N_A_893_101#_c_667_n N_A_1297_290#_c_845_n 4.06473e-19 $X=6.37 $Y=1.165
+ $X2=0 $Y2=0
cc_570 N_A_893_101#_c_673_n N_A_1297_290#_c_845_n 0.00957688f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_571 N_A_893_101#_c_673_n N_A_1297_290#_c_880_n 0.0070916f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_572 N_A_893_101#_c_667_n N_A_1297_290#_c_846_n 0.00621684f $X=6.37 $Y=1.165
+ $X2=0 $Y2=0
cc_573 N_A_893_101#_c_671_n N_A_1297_290#_c_846_n 0.00813837f $X=6.005 $Y=1.49
+ $X2=0 $Y2=0
cc_574 N_A_893_101#_c_673_n N_A_1297_290#_c_846_n 0.00695302f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_575 N_A_893_101#_c_673_n N_SET_B_M1026_g 0.00520105f $X=9.695 $Y=1.295 $X2=0
+ $Y2=0
cc_576 N_A_893_101#_c_673_n SET_B 0.0141171f $X=9.695 $Y=1.295 $X2=0 $Y2=0
cc_577 N_A_893_101#_c_681_n N_SET_B_c_1029_n 7.22754e-19 $X=9.74 $Y=2.455 $X2=0
+ $Y2=0
cc_578 N_A_893_101#_c_686_n N_SET_B_c_1029_n 0.0102124f $X=9.915 $Y=2.25 $X2=0
+ $Y2=0
cc_579 N_A_893_101#_c_675_n N_SET_B_c_1029_n 0.0114395f $X=9.84 $Y=1.295 $X2=0
+ $Y2=0
cc_580 N_A_893_101#_c_679_n N_SET_B_c_1029_n 0.0174461f $X=9.775 $Y=1.29 $X2=0
+ $Y2=0
cc_581 N_A_893_101#_c_673_n N_SET_B_c_1030_n 0.013249f $X=9.695 $Y=1.295 $X2=0
+ $Y2=0
cc_582 N_A_893_101#_c_673_n N_SET_B_c_1022_n 0.00489943f $X=9.695 $Y=1.295 $X2=0
+ $Y2=0
cc_583 N_A_893_101#_c_673_n N_SET_B_c_1034_n 0.00109848f $X=9.695 $Y=1.295 $X2=0
+ $Y2=0
cc_584 N_A_893_101#_c_673_n N_A_1216_457#_c_1154_n 0.00247074f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_585 N_A_893_101#_M1023_g N_A_1216_457#_c_1156_n 0.0189828f $X=6.515 $Y=0.445
+ $X2=0 $Y2=0
cc_586 N_A_893_101#_c_665_n N_A_1216_457#_c_1157_n 0.011075f $X=6.005 $Y=1.415
+ $X2=0 $Y2=0
cc_587 N_A_893_101#_c_667_n N_A_1216_457#_c_1157_n 0.00606684f $X=6.37 $Y=1.165
+ $X2=0 $Y2=0
cc_588 N_A_893_101#_c_673_n N_A_1216_457#_c_1157_n 0.0260853f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_589 N_A_893_101#_c_667_n N_A_1216_457#_c_1158_n 0.00368662f $X=6.37 $Y=1.165
+ $X2=0 $Y2=0
cc_590 N_A_893_101#_M1023_g N_A_1216_457#_c_1158_n 0.00616537f $X=6.515 $Y=0.445
+ $X2=0 $Y2=0
cc_591 N_A_893_101#_c_673_n N_A_1216_457#_c_1158_n 0.0438818f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_592 N_A_893_101#_c_667_n N_A_1216_457#_c_1159_n 0.0146868f $X=6.37 $Y=1.165
+ $X2=0 $Y2=0
cc_593 N_A_893_101#_M1023_g N_A_1216_457#_c_1159_n 7.66956e-19 $X=6.515 $Y=0.445
+ $X2=0 $Y2=0
cc_594 N_A_893_101#_c_673_n N_A_1216_457#_c_1159_n 0.00843506f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_595 N_A_893_101#_c_673_n N_A_1216_457#_c_1160_n 0.0249701f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_596 N_A_893_101#_c_673_n N_A_1650_21#_M1046_g 0.00135442f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_597 N_A_893_101#_c_673_n N_A_1650_21#_c_1253_n 0.0225201f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_598 N_A_893_101#_c_673_n N_A_1650_21#_c_1254_n 0.00978233f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_599 N_A_893_101#_M1018_g N_A_1650_21#_c_1255_n 7.94572e-19 $X=9.745 $Y=0.605
+ $X2=0 $Y2=0
cc_600 N_A_893_101#_c_673_n N_A_1650_21#_c_1255_n 0.021481f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_601 N_A_893_101#_M1018_g N_A_1650_21#_c_1257_n 0.0143861f $X=9.745 $Y=0.605
+ $X2=0 $Y2=0
cc_602 N_A_893_101#_c_672_n N_A_755_106#_c_1421_n 0.0187993f $X=4.61 $Y=0.78
+ $X2=0 $Y2=0
cc_603 N_A_893_101#_c_672_n N_A_755_106#_c_1423_n 0.0026033f $X=4.61 $Y=0.78
+ $X2=0 $Y2=0
cc_604 N_A_893_101#_c_664_n N_A_755_106#_M1042_g 0.0346282f $X=5.56 $Y=1.49
+ $X2=0 $Y2=0
cc_605 N_A_893_101#_c_672_n N_A_755_106#_M1042_g 0.010909f $X=4.61 $Y=0.78 $X2=0
+ $Y2=0
cc_606 N_A_893_101#_c_683_n N_A_755_106#_M1042_g 0.0199768f $X=4.7 $Y=2.43 $X2=0
+ $Y2=0
cc_607 N_A_893_101#_c_684_n N_A_755_106#_M1042_g 0.012635f $X=5.045 $Y=2 $X2=0
+ $Y2=0
cc_608 N_A_893_101#_c_685_n N_A_755_106#_M1042_g 0.00515835f $X=4.695 $Y=2 $X2=0
+ $Y2=0
cc_609 N_A_893_101#_c_674_n N_A_755_106#_M1042_g 0.004233f $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_610 N_A_893_101#_c_677_n N_A_755_106#_M1042_g 0.0110604f $X=5.395 $Y=1.58
+ $X2=0 $Y2=0
cc_611 N_A_893_101#_c_664_n N_A_755_106#_c_1425_n 0.0247611f $X=5.56 $Y=1.49
+ $X2=0 $Y2=0
cc_612 N_A_893_101#_c_667_n N_A_755_106#_c_1425_n 3.10308e-19 $X=6.37 $Y=1.165
+ $X2=0 $Y2=0
cc_613 N_A_893_101#_c_668_n N_A_755_106#_c_1425_n 0.00447088f $X=6.08 $Y=1.165
+ $X2=0 $Y2=0
cc_614 N_A_893_101#_c_673_n N_A_755_106#_c_1425_n 0.00665429f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_615 N_A_893_101#_c_677_n N_A_755_106#_c_1425_n 0.00693247f $X=5.395 $Y=1.58
+ $X2=0 $Y2=0
cc_616 N_A_893_101#_M1012_g N_A_755_106#_c_1436_n 0.00895007f $X=6.005 $Y=2.495
+ $X2=0 $Y2=0
cc_617 N_A_893_101#_c_663_n N_A_755_106#_c_1427_n 0.0041923f $X=5.93 $Y=1.49
+ $X2=0 $Y2=0
cc_618 N_A_893_101#_c_668_n N_A_755_106#_c_1427_n 0.0170286f $X=6.08 $Y=1.165
+ $X2=0 $Y2=0
cc_619 N_A_893_101#_c_673_n N_A_755_106#_c_1427_n 8.97469e-19 $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_620 N_A_893_101#_M1023_g N_A_755_106#_c_1429_n 0.0186678f $X=6.515 $Y=0.445
+ $X2=0 $Y2=0
cc_621 N_A_893_101#_M1012_g N_A_755_106#_M1043_g 0.0118797f $X=6.005 $Y=2.495
+ $X2=0 $Y2=0
cc_622 N_A_893_101#_c_681_n N_A_755_106#_c_1439_n 0.0107105f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_623 N_A_893_101#_c_681_n N_A_755_106#_M1035_g 0.015557f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_624 N_A_893_101#_c_686_n N_A_755_106#_M1035_g 0.00634664f $X=9.915 $Y=2.25
+ $X2=0 $Y2=0
cc_625 N_A_893_101#_c_679_n N_A_755_106#_M1035_g 2.54856e-19 $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_626 N_A_893_101#_c_681_n N_A_755_106#_c_1441_n 0.0197318f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_627 N_A_893_101#_c_686_n N_A_755_106#_c_1441_n 9.86368e-19 $X=9.915 $Y=2.25
+ $X2=0 $Y2=0
cc_628 N_A_893_101#_c_675_n N_A_755_106#_c_1441_n 4.25061e-19 $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_629 N_A_893_101#_c_678_n N_A_755_106#_c_1441_n 0.0181155f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_630 N_A_893_101#_c_679_n N_A_755_106#_c_1441_n 0.0177729f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_631 N_A_893_101#_c_673_n N_A_755_106#_c_1442_n 0.00466784f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_632 N_A_893_101#_c_679_n N_A_755_106#_c_1442_n 0.0051765f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_633 N_A_893_101#_M1018_g N_A_755_106#_M1027_g 0.0182003f $X=9.745 $Y=0.605
+ $X2=0 $Y2=0
cc_634 N_A_893_101#_c_678_n N_A_755_106#_M1027_g 0.0180735f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_635 N_A_893_101#_c_679_n N_A_755_106#_M1027_g 0.00468666f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_636 N_A_893_101#_c_672_n N_A_755_106#_c_1432_n 0.095109f $X=4.61 $Y=0.78
+ $X2=0 $Y2=0
cc_637 N_A_893_101#_c_672_n N_A_755_106#_c_1433_n 0.00480458f $X=4.61 $Y=0.78
+ $X2=0 $Y2=0
cc_638 N_A_893_101#_c_683_n N_A_755_106#_c_1446_n 0.0682329f $X=4.7 $Y=2.43
+ $X2=0 $Y2=0
cc_639 N_A_893_101#_c_685_n N_A_755_106#_c_1446_n 0.0143087f $X=4.695 $Y=2 $X2=0
+ $Y2=0
cc_640 N_A_893_101#_c_681_n N_A_2064_453#_M1017_g 0.0162468f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_641 N_A_893_101#_c_681_n N_A_2064_453#_c_1596_n 0.0137112f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_642 N_A_893_101#_c_681_n N_A_1861_431#_c_1765_n 0.0182033f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_643 N_A_893_101#_c_686_n N_A_1861_431#_c_1765_n 0.0272705f $X=9.915 $Y=2.25
+ $X2=0 $Y2=0
cc_644 N_A_893_101#_M1018_g N_A_1861_431#_c_1754_n 0.00433857f $X=9.745 $Y=0.605
+ $X2=0 $Y2=0
cc_645 N_A_893_101#_c_675_n N_A_1861_431#_c_1754_n 0.00256594f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_646 N_A_893_101#_c_678_n N_A_1861_431#_c_1754_n 8.80101e-19 $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_647 N_A_893_101#_c_679_n N_A_1861_431#_c_1754_n 0.0116137f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_648 N_A_893_101#_M1018_g N_A_1861_431#_c_1755_n 0.00322797f $X=9.745 $Y=0.605
+ $X2=0 $Y2=0
cc_649 N_A_893_101#_c_675_n N_A_1861_431#_c_1755_n 0.00558999f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_650 N_A_893_101#_c_678_n N_A_1861_431#_c_1755_n 6.62895e-19 $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_651 N_A_893_101#_c_679_n N_A_1861_431#_c_1755_n 0.0147898f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_652 N_A_893_101#_c_681_n N_A_1861_431#_c_1756_n 0.00572664f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_653 N_A_893_101#_c_686_n N_A_1861_431#_c_1756_n 0.0240749f $X=9.915 $Y=2.25
+ $X2=0 $Y2=0
cc_654 N_A_893_101#_c_679_n N_A_1861_431#_c_1756_n 0.0291318f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_655 N_A_893_101#_c_681_n N_A_1861_431#_c_1764_n 0.00174815f $X=9.74 $Y=2.455
+ $X2=0 $Y2=0
cc_656 N_A_893_101#_c_675_n N_A_1861_431#_c_1759_n 0.00189735f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_657 N_A_893_101#_c_678_n N_A_1861_431#_c_1759_n 4.00666e-19 $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_658 N_A_893_101#_c_679_n N_A_1861_431#_c_1759_n 0.0135405f $X=9.775 $Y=1.29
+ $X2=0 $Y2=0
cc_659 N_A_893_101#_M1012_g N_VPWR_c_2015_n 0.00371345f $X=6.005 $Y=2.495 $X2=0
+ $Y2=0
cc_660 N_A_893_101#_c_683_n N_VPWR_c_2015_n 0.0260022f $X=4.7 $Y=2.43 $X2=0
+ $Y2=0
cc_661 N_A_893_101#_c_676_n N_VPWR_c_2015_n 0.00111929f $X=5.395 $Y=1.58 $X2=0
+ $Y2=0
cc_662 N_A_893_101#_c_677_n N_VPWR_c_2015_n 0.0288289f $X=5.395 $Y=1.58 $X2=0
+ $Y2=0
cc_663 N_A_893_101#_c_683_n N_VPWR_c_2022_n 0.0131516f $X=4.7 $Y=2.43 $X2=0
+ $Y2=0
cc_664 N_A_893_101#_c_681_n N_VPWR_c_2032_n 0.00340772f $X=9.74 $Y=2.455 $X2=0
+ $Y2=0
cc_665 N_A_893_101#_M1012_g N_VPWR_c_2010_n 9.49986e-19 $X=6.005 $Y=2.495 $X2=0
+ $Y2=0
cc_666 N_A_893_101#_c_681_n N_VPWR_c_2010_n 0.00481437f $X=9.74 $Y=2.455 $X2=0
+ $Y2=0
cc_667 N_A_893_101#_c_683_n N_VPWR_c_2010_n 0.0120991f $X=4.7 $Y=2.43 $X2=0
+ $Y2=0
cc_668 N_A_893_101#_c_672_n N_A_204_119#_c_2210_n 0.0123913f $X=4.61 $Y=0.78
+ $X2=0 $Y2=0
cc_669 N_A_893_101#_c_663_n N_A_204_119#_c_2212_n 0.00102984f $X=5.93 $Y=1.49
+ $X2=0 $Y2=0
cc_670 N_A_893_101#_c_664_n N_A_204_119#_c_2212_n 4.20259e-19 $X=5.56 $Y=1.49
+ $X2=0 $Y2=0
cc_671 N_A_893_101#_c_673_n N_A_204_119#_c_2212_n 0.015236f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_672 N_A_893_101#_c_674_n N_A_204_119#_c_2212_n 0.00105873f $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_673 N_A_893_101#_c_677_n N_A_204_119#_c_2212_n 0.0180344f $X=5.395 $Y=1.58
+ $X2=0 $Y2=0
cc_674 N_A_893_101#_c_672_n N_A_204_119#_c_2213_n 0.00952293f $X=4.61 $Y=0.78
+ $X2=0 $Y2=0
cc_675 N_A_893_101#_c_674_n N_A_204_119#_c_2213_n 0.00252036f $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_676 N_A_893_101#_c_677_n N_A_204_119#_c_2213_n 0.0081945f $X=5.395 $Y=1.58
+ $X2=0 $Y2=0
cc_677 N_A_893_101#_c_663_n N_A_204_119#_c_2221_n 0.00303541f $X=5.93 $Y=1.49
+ $X2=0 $Y2=0
cc_678 N_A_893_101#_M1012_g N_A_204_119#_c_2221_n 0.00650457f $X=6.005 $Y=2.495
+ $X2=0 $Y2=0
cc_679 N_A_893_101#_c_663_n N_A_204_119#_c_2216_n 0.00834547f $X=5.93 $Y=1.49
+ $X2=0 $Y2=0
cc_680 N_A_893_101#_c_665_n N_A_204_119#_c_2216_n 0.00440497f $X=6.005 $Y=1.415
+ $X2=0 $Y2=0
cc_681 N_A_893_101#_M1012_g N_A_204_119#_c_2216_n 0.0153849f $X=6.005 $Y=2.495
+ $X2=0 $Y2=0
cc_682 N_A_893_101#_c_668_n N_A_204_119#_c_2216_n 0.00424127f $X=6.08 $Y=1.165
+ $X2=0 $Y2=0
cc_683 N_A_893_101#_M1023_g N_A_204_119#_c_2216_n 2.26516e-19 $X=6.515 $Y=0.445
+ $X2=0 $Y2=0
cc_684 N_A_893_101#_c_671_n N_A_204_119#_c_2216_n 0.00160772f $X=6.005 $Y=1.49
+ $X2=0 $Y2=0
cc_685 N_A_893_101#_c_673_n N_A_204_119#_c_2216_n 0.0168655f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_686 N_A_893_101#_c_674_n N_A_204_119#_c_2216_n 5.43297e-19 $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_687 N_A_893_101#_c_676_n N_A_204_119#_c_2216_n 0.00183347f $X=5.395 $Y=1.58
+ $X2=0 $Y2=0
cc_688 N_A_893_101#_c_677_n N_A_204_119#_c_2216_n 0.047423f $X=5.395 $Y=1.58
+ $X2=0 $Y2=0
cc_689 N_A_893_101#_c_663_n N_A_204_119#_c_2217_n 0.00179456f $X=5.93 $Y=1.49
+ $X2=0 $Y2=0
cc_690 N_A_893_101#_M1023_g N_A_204_119#_c_2217_n 5.32524e-19 $X=6.515 $Y=0.445
+ $X2=0 $Y2=0
cc_691 N_A_893_101#_c_673_n N_A_204_119#_c_2217_n 0.00398953f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_692 N_A_893_101#_M1018_g N_VGND_c_2460_n 9.62076e-19 $X=9.745 $Y=0.605 $X2=0
+ $Y2=0
cc_693 N_A_893_101#_M1023_g N_VGND_c_2470_n 0.00549284f $X=6.515 $Y=0.445 $X2=0
+ $Y2=0
cc_694 N_A_893_101#_M1018_g N_VGND_c_2474_n 0.00327726f $X=9.745 $Y=0.605 $X2=0
+ $Y2=0
cc_695 N_A_893_101#_M1023_g N_VGND_c_2480_n 0.00995098f $X=6.515 $Y=0.445 $X2=0
+ $Y2=0
cc_696 N_A_893_101#_M1018_g N_VGND_c_2480_n 0.00577104f $X=9.745 $Y=0.605 $X2=0
+ $Y2=0
cc_697 N_A_893_101#_c_673_n N_A_1492_47#_c_2640_n 0.0010329f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_698 N_A_1297_290#_M1010_g N_SET_B_M1026_g 0.0347726f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_699 N_A_1297_290#_c_852_n N_SET_B_M1040_g 0.0144519f $X=7.465 $Y=2.415 $X2=0
+ $Y2=0
cc_700 N_A_1297_290#_c_866_n N_SET_B_M1040_g 0.00202937f $X=7.63 $Y=2.13 $X2=0
+ $Y2=0
cc_701 N_A_1297_290#_c_887_p N_SET_B_M1040_g 0.00406107f $X=7.63 $Y=2.33 $X2=0
+ $Y2=0
cc_702 N_A_1297_290#_c_846_n N_SET_B_M1040_g 0.0263468f $X=6.825 $Y=1.615 $X2=0
+ $Y2=0
cc_703 N_A_1297_290#_M1016_g N_SET_B_c_1027_n 0.00171885f $X=6.825 $Y=2.495
+ $X2=0 $Y2=0
cc_704 N_A_1297_290#_c_851_n N_SET_B_c_1027_n 0.00731172f $X=6.57 $Y=2.33 $X2=0
+ $Y2=0
cc_705 N_A_1297_290#_M1010_g SET_B 0.00340306f $X=6.875 $Y=0.445 $X2=0 $Y2=0
cc_706 N_A_1297_290#_c_851_n SET_B 4.24405e-19 $X=6.57 $Y=2.33 $X2=0 $Y2=0
cc_707 N_A_1297_290#_c_852_n SET_B 0.00357092f $X=7.465 $Y=2.415 $X2=0 $Y2=0
cc_708 N_A_1297_290#_c_866_n SET_B 0.00281255f $X=7.63 $Y=2.13 $X2=0 $Y2=0
cc_709 N_A_1297_290#_c_842_n SET_B 0.00268865f $X=8.26 $Y=1.96 $X2=0 $Y2=0
cc_710 N_A_1297_290#_c_845_n SET_B 0.0252769f $X=6.65 $Y=1.615 $X2=0 $Y2=0
cc_711 N_A_1297_290#_c_846_n SET_B 0.00168245f $X=6.825 $Y=1.615 $X2=0 $Y2=0
cc_712 N_A_1297_290#_c_852_n N_SET_B_c_1029_n 0.00833869f $X=7.465 $Y=2.415
+ $X2=0 $Y2=0
cc_713 N_A_1297_290#_c_866_n N_SET_B_c_1029_n 0.0341044f $X=7.63 $Y=2.13 $X2=0
+ $Y2=0
cc_714 N_A_1297_290#_c_867_n N_SET_B_c_1029_n 0.0310818f $X=8.175 $Y=2.045 $X2=0
+ $Y2=0
cc_715 N_A_1297_290#_c_854_n N_SET_B_c_1029_n 0.0819588f $X=9.03 $Y=2.045 $X2=0
+ $Y2=0
cc_716 N_A_1297_290#_c_844_n N_SET_B_c_1029_n 2.28044e-19 $X=9.195 $Y=1.29 $X2=0
+ $Y2=0
cc_717 N_A_1297_290#_c_903_p N_SET_B_c_1029_n 0.0189773f $X=8.26 $Y=2.045 $X2=0
+ $Y2=0
cc_718 N_A_1297_290#_M1016_g N_SET_B_c_1030_n 0.00429414f $X=6.825 $Y=2.495
+ $X2=0 $Y2=0
cc_719 N_A_1297_290#_c_851_n N_SET_B_c_1030_n 0.00656879f $X=6.57 $Y=2.33 $X2=0
+ $Y2=0
cc_720 N_A_1297_290#_c_852_n N_SET_B_c_1030_n 0.00806122f $X=7.465 $Y=2.415
+ $X2=0 $Y2=0
cc_721 N_A_1297_290#_c_846_n N_SET_B_c_1030_n 9.72579e-19 $X=6.825 $Y=1.615
+ $X2=0 $Y2=0
cc_722 N_A_1297_290#_M1010_g N_SET_B_c_1022_n 0.0138548f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_723 N_A_1297_290#_c_852_n N_SET_B_c_1022_n 6.59835e-19 $X=7.465 $Y=2.415
+ $X2=0 $Y2=0
cc_724 N_A_1297_290#_c_845_n N_SET_B_c_1022_n 2.01141e-19 $X=6.65 $Y=1.615 $X2=0
+ $Y2=0
cc_725 N_A_1297_290#_c_846_n N_SET_B_c_1022_n 0.0050108f $X=6.825 $Y=1.615 $X2=0
+ $Y2=0
cc_726 N_A_1297_290#_M1016_g N_SET_B_c_1034_n 0.00615414f $X=6.825 $Y=2.495
+ $X2=0 $Y2=0
cc_727 N_A_1297_290#_c_851_n N_SET_B_c_1034_n 0.0110845f $X=6.57 $Y=2.33 $X2=0
+ $Y2=0
cc_728 N_A_1297_290#_c_852_n N_SET_B_c_1034_n 0.0177472f $X=7.465 $Y=2.415 $X2=0
+ $Y2=0
cc_729 N_A_1297_290#_c_866_n N_SET_B_c_1034_n 0.00648569f $X=7.63 $Y=2.13 $X2=0
+ $Y2=0
cc_730 N_A_1297_290#_c_887_p N_SET_B_c_1034_n 8.06547e-19 $X=7.63 $Y=2.33 $X2=0
+ $Y2=0
cc_731 N_A_1297_290#_c_846_n N_SET_B_c_1034_n 0.00150474f $X=6.825 $Y=1.615
+ $X2=0 $Y2=0
cc_732 N_A_1297_290#_c_842_n N_A_1216_457#_M1001_g 0.00357776f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_733 N_A_1297_290#_c_852_n N_A_1216_457#_M1024_g 0.00831339f $X=7.465 $Y=2.415
+ $X2=0 $Y2=0
cc_734 N_A_1297_290#_c_866_n N_A_1216_457#_M1024_g 8.23351e-19 $X=7.63 $Y=2.13
+ $X2=0 $Y2=0
cc_735 N_A_1297_290#_c_887_p N_A_1216_457#_M1024_g 0.00385909f $X=7.63 $Y=2.33
+ $X2=0 $Y2=0
cc_736 N_A_1297_290#_c_867_n N_A_1216_457#_M1024_g 0.0118227f $X=8.175 $Y=2.045
+ $X2=0 $Y2=0
cc_737 N_A_1297_290#_c_842_n N_A_1216_457#_M1024_g 0.00421769f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_738 N_A_1297_290#_c_866_n N_A_1216_457#_c_1155_n 5.19222e-19 $X=7.63 $Y=2.13
+ $X2=0 $Y2=0
cc_739 N_A_1297_290#_c_867_n N_A_1216_457#_c_1155_n 0.00165163f $X=8.175
+ $Y=2.045 $X2=0 $Y2=0
cc_740 N_A_1297_290#_M1010_g N_A_1216_457#_c_1156_n 0.0025485f $X=6.875 $Y=0.445
+ $X2=0 $Y2=0
cc_741 N_A_1297_290#_M1016_g N_A_1216_457#_c_1157_n 5.20892e-19 $X=6.825
+ $Y=2.495 $X2=0 $Y2=0
cc_742 N_A_1297_290#_M1010_g N_A_1216_457#_c_1157_n 0.00290364f $X=6.875
+ $Y=0.445 $X2=0 $Y2=0
cc_743 N_A_1297_290#_c_851_n N_A_1216_457#_c_1157_n 0.037443f $X=6.57 $Y=2.33
+ $X2=0 $Y2=0
cc_744 N_A_1297_290#_c_845_n N_A_1216_457#_c_1157_n 0.0229991f $X=6.65 $Y=1.615
+ $X2=0 $Y2=0
cc_745 N_A_1297_290#_c_846_n N_A_1216_457#_c_1157_n 0.00122188f $X=6.825
+ $Y=1.615 $X2=0 $Y2=0
cc_746 N_A_1297_290#_M1010_g N_A_1216_457#_c_1158_n 0.0150166f $X=6.875 $Y=0.445
+ $X2=0 $Y2=0
cc_747 N_A_1297_290#_c_845_n N_A_1216_457#_c_1158_n 0.0113441f $X=6.65 $Y=1.615
+ $X2=0 $Y2=0
cc_748 N_A_1297_290#_c_846_n N_A_1216_457#_c_1158_n 0.00499015f $X=6.825
+ $Y=1.615 $X2=0 $Y2=0
cc_749 N_A_1297_290#_c_866_n N_A_1216_457#_c_1160_n 0.00266411f $X=7.63 $Y=2.13
+ $X2=0 $Y2=0
cc_750 N_A_1297_290#_c_867_n N_A_1216_457#_c_1160_n 0.00705511f $X=8.175
+ $Y=2.045 $X2=0 $Y2=0
cc_751 N_A_1297_290#_c_842_n N_A_1216_457#_c_1160_n 0.0475041f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_752 N_A_1297_290#_c_880_n N_A_1216_457#_c_1160_n 0.00304572f $X=8.26 $Y=0.73
+ $X2=0 $Y2=0
cc_753 N_A_1297_290#_c_842_n N_A_1216_457#_c_1161_n 0.00369466f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_754 N_A_1297_290#_c_880_n N_A_1216_457#_c_1161_n 0.00170657f $X=8.26 $Y=0.73
+ $X2=0 $Y2=0
cc_755 N_A_1297_290#_c_842_n N_A_1650_21#_c_1248_n 0.0036908f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_756 N_A_1297_290#_c_880_n N_A_1650_21#_c_1248_n 0.00865968f $X=8.26 $Y=0.73
+ $X2=0 $Y2=0
cc_757 N_A_1297_290#_c_840_n N_A_1650_21#_M1046_g 0.0418048f $X=8.83 $Y=1.6
+ $X2=0 $Y2=0
cc_758 N_A_1297_290#_c_852_n N_A_1650_21#_M1046_g 0.00120132f $X=7.465 $Y=2.415
+ $X2=0 $Y2=0
cc_759 N_A_1297_290#_c_887_p N_A_1650_21#_M1046_g 9.16241e-19 $X=7.63 $Y=2.33
+ $X2=0 $Y2=0
cc_760 N_A_1297_290#_c_842_n N_A_1650_21#_M1046_g 0.018591f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_761 N_A_1297_290#_c_854_n N_A_1650_21#_M1046_g 0.00577775f $X=9.03 $Y=2.045
+ $X2=0 $Y2=0
cc_762 N_A_1297_290#_c_843_n N_A_1650_21#_M1046_g 0.00157368f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_763 N_A_1297_290#_c_844_n N_A_1650_21#_M1046_g 0.00333592f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_764 N_A_1297_290#_c_903_p N_A_1650_21#_M1046_g 0.00866526f $X=8.26 $Y=2.045
+ $X2=0 $Y2=0
cc_765 N_A_1297_290#_c_840_n N_A_1650_21#_c_1253_n 9.83524e-19 $X=8.83 $Y=1.6
+ $X2=0 $Y2=0
cc_766 N_A_1297_290#_M1008_g N_A_1650_21#_c_1253_n 0.00188239f $X=9.325 $Y=0.605
+ $X2=0 $Y2=0
cc_767 N_A_1297_290#_c_842_n N_A_1650_21#_c_1253_n 0.0245129f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_768 N_A_1297_290#_c_854_n N_A_1650_21#_c_1253_n 0.00291753f $X=9.03 $Y=2.045
+ $X2=0 $Y2=0
cc_769 N_A_1297_290#_c_843_n N_A_1650_21#_c_1253_n 0.0109261f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_770 N_A_1297_290#_c_844_n N_A_1650_21#_c_1253_n 6.60849e-19 $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_771 N_A_1297_290#_c_840_n N_A_1650_21#_c_1254_n 0.00935083f $X=8.83 $Y=1.6
+ $X2=0 $Y2=0
cc_772 N_A_1297_290#_M1008_g N_A_1650_21#_c_1254_n 0.00451692f $X=9.325 $Y=0.605
+ $X2=0 $Y2=0
cc_773 N_A_1297_290#_c_842_n N_A_1650_21#_c_1254_n 0.00839028f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_774 N_A_1297_290#_c_854_n N_A_1650_21#_c_1254_n 0.00222078f $X=9.03 $Y=2.045
+ $X2=0 $Y2=0
cc_775 N_A_1297_290#_c_843_n N_A_1650_21#_c_1254_n 7.02243e-19 $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_776 N_A_1297_290#_c_844_n N_A_1650_21#_c_1254_n 0.0128574f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_777 N_A_1297_290#_c_840_n N_A_1650_21#_c_1255_n 0.00470759f $X=8.83 $Y=1.6
+ $X2=0 $Y2=0
cc_778 N_A_1297_290#_M1008_g N_A_1650_21#_c_1255_n 0.0132197f $X=9.325 $Y=0.605
+ $X2=0 $Y2=0
cc_779 N_A_1297_290#_c_843_n N_A_1650_21#_c_1255_n 0.0228484f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_780 N_A_1297_290#_c_844_n N_A_1650_21#_c_1255_n 0.00151583f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_781 N_A_1297_290#_c_842_n N_A_1650_21#_c_1256_n 0.0099412f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_782 N_A_1297_290#_c_880_n N_A_1650_21#_c_1256_n 0.00313763f $X=8.26 $Y=0.73
+ $X2=0 $Y2=0
cc_783 N_A_1297_290#_M1008_g N_A_1650_21#_c_1258_n 7.8785e-19 $X=9.325 $Y=0.605
+ $X2=0 $Y2=0
cc_784 N_A_1297_290#_M1016_g N_A_755_106#_M1043_g 0.0358479f $X=6.825 $Y=2.495
+ $X2=0 $Y2=0
cc_785 N_A_1297_290#_c_851_n N_A_755_106#_M1043_g 0.00327053f $X=6.57 $Y=2.33
+ $X2=0 $Y2=0
cc_786 N_A_1297_290#_c_972_p N_A_755_106#_M1043_g 0.00418265f $X=6.655 $Y=2.415
+ $X2=0 $Y2=0
cc_787 N_A_1297_290#_c_846_n N_A_755_106#_M1043_g 7.85634e-19 $X=6.825 $Y=1.615
+ $X2=0 $Y2=0
cc_788 N_A_1297_290#_M1016_g N_A_755_106#_c_1439_n 0.00861299f $X=6.825 $Y=2.495
+ $X2=0 $Y2=0
cc_789 N_A_1297_290#_M1031_g N_A_755_106#_c_1439_n 0.00894529f $X=8.755 $Y=2.285
+ $X2=0 $Y2=0
cc_790 N_A_1297_290#_c_852_n N_A_755_106#_c_1439_n 0.00915571f $X=7.465 $Y=2.415
+ $X2=0 $Y2=0
cc_791 N_A_1297_290#_c_972_p N_A_755_106#_c_1439_n 0.00146735f $X=6.655 $Y=2.415
+ $X2=0 $Y2=0
cc_792 N_A_1297_290#_c_854_n N_A_755_106#_M1035_g 0.00954352f $X=9.03 $Y=2.045
+ $X2=0 $Y2=0
cc_793 N_A_1297_290#_M1031_g N_A_755_106#_c_1442_n 0.0380542f $X=8.755 $Y=2.285
+ $X2=0 $Y2=0
cc_794 N_A_1297_290#_c_854_n N_A_755_106#_c_1442_n 0.00510349f $X=9.03 $Y=2.045
+ $X2=0 $Y2=0
cc_795 N_A_1297_290#_c_843_n N_A_755_106#_c_1442_n 0.0083207f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_796 N_A_1297_290#_c_844_n N_A_755_106#_c_1442_n 0.00699541f $X=9.195 $Y=1.29
+ $X2=0 $Y2=0
cc_797 N_A_1297_290#_M1031_g N_A_1861_431#_c_1764_n 7.28369e-19 $X=8.755
+ $Y=2.285 $X2=0 $Y2=0
cc_798 N_A_1297_290#_c_854_n N_A_1861_431#_c_1764_n 0.00195818f $X=9.03 $Y=2.045
+ $X2=0 $Y2=0
cc_799 N_A_1297_290#_c_852_n N_VPWR_M1016_d 0.00761269f $X=7.465 $Y=2.415 $X2=0
+ $Y2=0
cc_800 N_A_1297_290#_c_854_n N_VPWR_M1046_d 0.00410544f $X=9.03 $Y=2.045 $X2=0
+ $Y2=0
cc_801 N_A_1297_290#_M1016_g N_VPWR_c_2016_n 0.00366822f $X=6.825 $Y=2.495 $X2=0
+ $Y2=0
cc_802 N_A_1297_290#_c_852_n N_VPWR_c_2016_n 0.0261733f $X=7.465 $Y=2.415 $X2=0
+ $Y2=0
cc_803 N_A_1297_290#_M1031_g N_VPWR_c_2017_n 0.0120439f $X=8.755 $Y=2.285 $X2=0
+ $Y2=0
cc_804 N_A_1297_290#_c_852_n N_VPWR_c_2017_n 0.0110626f $X=7.465 $Y=2.415 $X2=0
+ $Y2=0
cc_805 N_A_1297_290#_c_887_p N_VPWR_c_2017_n 5.31704e-19 $X=7.63 $Y=2.33 $X2=0
+ $Y2=0
cc_806 N_A_1297_290#_c_854_n N_VPWR_c_2017_n 0.0146903f $X=9.03 $Y=2.045 $X2=0
+ $Y2=0
cc_807 N_A_1297_290#_c_852_n N_VPWR_c_2031_n 0.00699294f $X=7.465 $Y=2.415 $X2=0
+ $Y2=0
cc_808 N_A_1297_290#_M1016_g N_VPWR_c_2010_n 9.49986e-19 $X=6.825 $Y=2.495 $X2=0
+ $Y2=0
cc_809 N_A_1297_290#_M1031_g N_VPWR_c_2010_n 7.97988e-19 $X=8.755 $Y=2.285 $X2=0
+ $Y2=0
cc_810 N_A_1297_290#_c_852_n N_VPWR_c_2010_n 0.0239816f $X=7.465 $Y=2.415 $X2=0
+ $Y2=0
cc_811 N_A_1297_290#_c_972_p N_VPWR_c_2010_n 0.00596597f $X=6.655 $Y=2.415 $X2=0
+ $Y2=0
cc_812 N_A_1297_290#_c_851_n A_1302_457# 4.89857e-19 $X=6.57 $Y=2.33 $X2=-0.19
+ $Y2=-0.245
cc_813 N_A_1297_290#_c_852_n A_1302_457# 8.81966e-19 $X=7.465 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_814 N_A_1297_290#_c_972_p A_1302_457# 0.00132393f $X=6.655 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_815 N_A_1297_290#_c_867_n A_1584_373# 0.0108213f $X=8.175 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_816 N_A_1297_290#_c_842_n A_1584_373# 0.00116286f $X=8.26 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_817 N_A_1297_290#_c_903_p A_1584_373# 7.66879e-19 $X=8.26 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_818 N_A_1297_290#_c_854_n A_1766_373# 0.00857814f $X=9.03 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_819 N_A_1297_290#_c_843_n A_1766_373# 0.0012063f $X=9.195 $Y=1.29 $X2=-0.19
+ $Y2=-0.245
cc_820 N_A_1297_290#_M1010_g N_VGND_c_2459_n 0.00767498f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_821 N_A_1297_290#_M1008_g N_VGND_c_2460_n 0.00846366f $X=9.325 $Y=0.605 $X2=0
+ $Y2=0
cc_822 N_A_1297_290#_M1010_g N_VGND_c_2470_n 0.00585385f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_823 N_A_1297_290#_M1008_g N_VGND_c_2474_n 0.0048079f $X=9.325 $Y=0.605 $X2=0
+ $Y2=0
cc_824 N_A_1297_290#_M1001_d N_VGND_c_2480_n 0.00289884f $X=7.89 $Y=0.235 $X2=0
+ $Y2=0
cc_825 N_A_1297_290#_M1010_g N_VGND_c_2480_n 0.0109146f $X=6.875 $Y=0.445 $X2=0
+ $Y2=0
cc_826 N_A_1297_290#_M1008_g N_VGND_c_2480_n 0.00454109f $X=9.325 $Y=0.605 $X2=0
+ $Y2=0
cc_827 N_A_1297_290#_c_842_n N_A_1492_47#_c_2640_n 0.00112274f $X=8.26 $Y=1.96
+ $X2=0 $Y2=0
cc_828 N_A_1297_290#_M1001_d N_A_1492_47#_c_2639_n 0.0049838f $X=7.89 $Y=0.235
+ $X2=0 $Y2=0
cc_829 N_A_1297_290#_M1008_g N_A_1492_47#_c_2639_n 4.44372e-19 $X=9.325 $Y=0.605
+ $X2=0 $Y2=0
cc_830 N_A_1297_290#_c_880_n N_A_1492_47#_c_2639_n 0.0222108f $X=8.26 $Y=0.73
+ $X2=0 $Y2=0
cc_831 N_SET_B_M1026_g N_A_1216_457#_M1001_g 0.0256445f $X=7.385 $Y=0.555 $X2=0
+ $Y2=0
cc_832 SET_B N_A_1216_457#_M1024_g 9.04246e-19 $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_833 N_SET_B_c_1022_n N_A_1216_457#_M1024_g 0.0181697f $X=7.325 $Y=1.54 $X2=0
+ $Y2=0
cc_834 SET_B N_A_1216_457#_c_1154_n 0.0019178f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_835 N_SET_B_c_1022_n N_A_1216_457#_c_1154_n 0.0199981f $X=7.325 $Y=1.54 $X2=0
+ $Y2=0
cc_836 N_SET_B_M1026_g N_A_1216_457#_c_1158_n 0.0143784f $X=7.385 $Y=0.555 $X2=0
+ $Y2=0
cc_837 SET_B N_A_1216_457#_c_1158_n 0.0295012f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_838 N_SET_B_c_1022_n N_A_1216_457#_c_1158_n 0.00412671f $X=7.325 $Y=1.54
+ $X2=0 $Y2=0
cc_839 N_SET_B_M1026_g N_A_1216_457#_c_1160_n 0.00168376f $X=7.385 $Y=0.555
+ $X2=0 $Y2=0
cc_840 SET_B N_A_1216_457#_c_1160_n 0.024983f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_841 N_SET_B_c_1029_n N_A_1216_457#_c_1160_n 0.00220202f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_842 N_SET_B_c_1022_n N_A_1216_457#_c_1160_n 3.691e-19 $X=7.325 $Y=1.54 $X2=0
+ $Y2=0
cc_843 N_SET_B_M1026_g N_A_1216_457#_c_1161_n 0.0199641f $X=7.385 $Y=0.555 $X2=0
+ $Y2=0
cc_844 N_SET_B_M1011_g N_A_1650_21#_c_1259_n 9.38995e-19 $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_845 N_SET_B_M1011_g N_A_1650_21#_c_1260_n 0.015f $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_846 N_SET_B_M1011_g N_A_1650_21#_c_1266_n 0.00358112f $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_847 N_SET_B_M1040_g N_A_755_106#_c_1439_n 0.00856127f $X=7.415 $Y=2.285 $X2=0
+ $Y2=0
cc_848 N_SET_B_c_1029_n N_A_755_106#_c_1441_n 0.00642817f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_849 N_SET_B_c_1029_n N_A_755_106#_c_1442_n 0.0091984f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_850 N_SET_B_M1011_g N_A_2064_453#_M1009_g 0.0278312f $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_851 N_SET_B_M1020_g N_A_2064_453#_c_1596_n 0.00867142f $X=11.39 $Y=2.675
+ $X2=0 $Y2=0
cc_852 N_SET_B_c_1029_n N_A_2064_453#_c_1596_n 0.00823157f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_853 N_SET_B_c_1033_n N_A_2064_453#_c_1596_n 4.38352e-19 $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_854 N_SET_B_c_1019_n N_A_2064_453#_c_1597_n 0.00113999f $X=11.39 $Y=2.095
+ $X2=0 $Y2=0
cc_855 N_SET_B_M1020_g N_A_2064_453#_c_1597_n 0.00105241f $X=11.39 $Y=2.675
+ $X2=0 $Y2=0
cc_856 N_SET_B_c_1029_n N_A_2064_453#_c_1597_n 0.026261f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_857 N_SET_B_c_1021_n N_A_2064_453#_c_1597_n 5.61248e-19 $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_858 N_SET_B_c_1033_n N_A_2064_453#_c_1597_n 0.0222027f $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_859 N_SET_B_M1011_g N_A_2064_453#_c_1598_n 6.92146e-19 $X=11.32 $Y=0.605
+ $X2=0 $Y2=0
cc_860 N_SET_B_c_1019_n N_A_2064_453#_c_1598_n 0.0214129f $X=11.39 $Y=2.095
+ $X2=0 $Y2=0
cc_861 N_SET_B_c_1033_n N_A_2064_453#_c_1598_n 0.00113205f $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_862 N_SET_B_c_1019_n N_A_2064_453#_c_1599_n 0.00128788f $X=11.39 $Y=2.095
+ $X2=0 $Y2=0
cc_863 N_SET_B_M1020_g N_A_2064_453#_c_1599_n 0.0146269f $X=11.39 $Y=2.675 $X2=0
+ $Y2=0
cc_864 N_SET_B_c_1029_n N_A_2064_453#_c_1599_n 0.00941347f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_865 N_SET_B_c_1021_n N_A_2064_453#_c_1599_n 0.00266617f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_866 N_SET_B_c_1033_n N_A_2064_453#_c_1599_n 0.0187219f $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_867 N_SET_B_M1011_g N_A_1861_431#_M1028_g 0.0554858f $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_868 N_SET_B_c_1019_n N_A_1861_431#_M1021_g 0.0246832f $X=11.39 $Y=2.095 $X2=0
+ $Y2=0
cc_869 N_SET_B_c_1021_n N_A_1861_431#_M1021_g 5.25533e-19 $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_870 N_SET_B_c_1033_n N_A_1861_431#_M1021_g 9.25383e-19 $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_871 N_SET_B_c_1029_n N_A_1861_431#_c_1765_n 0.00761205f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_872 N_SET_B_c_1029_n N_A_1861_431#_c_1756_n 0.0191512f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_873 N_SET_B_M1011_g N_A_1861_431#_c_1757_n 0.0119301f $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_874 N_SET_B_c_1019_n N_A_1861_431#_c_1757_n 0.00278395f $X=11.39 $Y=2.095
+ $X2=0 $Y2=0
cc_875 N_SET_B_c_1029_n N_A_1861_431#_c_1757_n 0.0150984f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_876 N_SET_B_c_1021_n N_A_1861_431#_c_1757_n 0.00196756f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_877 N_SET_B_c_1033_n N_A_1861_431#_c_1757_n 0.0166893f $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_878 N_SET_B_M1011_g N_A_1861_431#_c_1758_n 0.0038948f $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_879 N_SET_B_c_1029_n N_A_1861_431#_c_1764_n 0.00968673f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_880 N_SET_B_c_1029_n N_A_1861_431#_c_1759_n 0.00345536f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_881 N_SET_B_M1011_g N_A_1861_431#_c_1760_n 0.00115038f $X=11.32 $Y=0.605
+ $X2=0 $Y2=0
cc_882 N_SET_B_c_1019_n N_A_1861_431#_c_1760_n 0.00178491f $X=11.39 $Y=2.095
+ $X2=0 $Y2=0
cc_883 N_SET_B_c_1021_n N_A_1861_431#_c_1760_n 0.00362507f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_884 N_SET_B_c_1033_n N_A_1861_431#_c_1760_n 0.0197887f $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_885 N_SET_B_c_1019_n N_A_1861_431#_c_1761_n 0.0147738f $X=11.39 $Y=2.095
+ $X2=0 $Y2=0
cc_886 N_SET_B_c_1033_n N_A_1861_431#_c_1761_n 3.59459e-19 $X=11.245 $Y=1.93
+ $X2=0 $Y2=0
cc_887 N_SET_B_c_1027_n N_VPWR_M1016_d 0.00229658f $X=7.08 $Y=1.95 $X2=0 $Y2=0
cc_888 N_SET_B_c_1029_n N_VPWR_M1016_d 0.00287448f $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_889 N_SET_B_c_1030_n N_VPWR_M1016_d 0.00139146f $X=7.105 $Y=2.035 $X2=0 $Y2=0
cc_890 N_SET_B_c_1034_n N_VPWR_M1016_d 0.004476f $X=7.08 $Y=2.05 $X2=0 $Y2=0
cc_891 N_SET_B_M1040_g N_VPWR_c_2016_n 0.00354178f $X=7.415 $Y=2.285 $X2=0 $Y2=0
cc_892 N_SET_B_c_1029_n N_VPWR_c_2017_n 0.00264269f $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_893 N_SET_B_M1020_g N_VPWR_c_2018_n 0.0113596f $X=11.39 $Y=2.675 $X2=0 $Y2=0
cc_894 N_SET_B_M1020_g N_VPWR_c_2024_n 0.00486043f $X=11.39 $Y=2.675 $X2=0 $Y2=0
cc_895 N_SET_B_M1040_g N_VPWR_c_2010_n 9.49986e-19 $X=7.415 $Y=2.285 $X2=0 $Y2=0
cc_896 N_SET_B_M1020_g N_VPWR_c_2010_n 0.00482043f $X=11.39 $Y=2.675 $X2=0 $Y2=0
cc_897 N_SET_B_M1026_g N_VGND_c_2459_n 0.00408627f $X=7.385 $Y=0.555 $X2=0 $Y2=0
cc_898 N_SET_B_M1011_g N_VGND_c_2461_n 0.00929942f $X=11.32 $Y=0.605 $X2=0 $Y2=0
cc_899 N_SET_B_M1026_g N_VGND_c_2472_n 0.0054778f $X=7.385 $Y=0.555 $X2=0 $Y2=0
cc_900 N_SET_B_M1011_g N_VGND_c_2478_n 0.00502664f $X=11.32 $Y=0.605 $X2=0 $Y2=0
cc_901 N_SET_B_M1026_g N_VGND_c_2480_n 0.0101836f $X=7.385 $Y=0.555 $X2=0 $Y2=0
cc_902 N_SET_B_M1011_g N_VGND_c_2480_n 0.0103357f $X=11.32 $Y=0.605 $X2=0 $Y2=0
cc_903 N_SET_B_M1026_g N_A_1492_47#_c_2640_n 0.00543609f $X=7.385 $Y=0.555 $X2=0
+ $Y2=0
cc_904 N_SET_B_M1026_g N_A_1492_47#_c_2646_n 0.00343647f $X=7.385 $Y=0.555 $X2=0
+ $Y2=0
cc_905 N_SET_B_M1011_g N_A_2279_57#_c_2670_n 0.00501801f $X=11.32 $Y=0.605 $X2=0
+ $Y2=0
cc_906 N_A_1216_457#_M1001_g N_A_1650_21#_c_1248_n 0.0245451f $X=7.815 $Y=0.555
+ $X2=0 $Y2=0
cc_907 N_A_1216_457#_M1024_g N_A_1650_21#_M1046_g 0.0399329f $X=7.845 $Y=2.285
+ $X2=0 $Y2=0
cc_908 N_A_1216_457#_c_1154_n N_A_1650_21#_M1046_g 0.0199878f $X=7.865 $Y=1.53
+ $X2=0 $Y2=0
cc_909 N_A_1216_457#_c_1160_n N_A_1650_21#_c_1254_n 5.92586e-19 $X=7.865 $Y=1.19
+ $X2=0 $Y2=0
cc_910 N_A_1216_457#_c_1161_n N_A_1650_21#_c_1254_n 0.0199878f $X=7.865 $Y=1.19
+ $X2=0 $Y2=0
cc_911 N_A_1216_457#_c_1157_n N_A_755_106#_c_1436_n 0.00265981f $X=6.22 $Y=2.495
+ $X2=0 $Y2=0
cc_912 N_A_1216_457#_c_1156_n N_A_755_106#_c_1426_n 5.37013e-19 $X=6.3 $Y=0.47
+ $X2=0 $Y2=0
cc_913 N_A_1216_457#_c_1156_n N_A_755_106#_c_1427_n 0.0045093f $X=6.3 $Y=0.47
+ $X2=0 $Y2=0
cc_914 N_A_1216_457#_c_1156_n N_A_755_106#_c_1429_n 0.00625553f $X=6.3 $Y=0.47
+ $X2=0 $Y2=0
cc_915 N_A_1216_457#_c_1157_n N_A_755_106#_M1043_g 0.00129909f $X=6.22 $Y=2.495
+ $X2=0 $Y2=0
cc_916 N_A_1216_457#_M1024_g N_A_755_106#_c_1439_n 0.00894493f $X=7.845 $Y=2.285
+ $X2=0 $Y2=0
cc_917 N_A_1216_457#_c_1157_n N_VPWR_c_2016_n 5.7929e-19 $X=6.22 $Y=2.495 $X2=0
+ $Y2=0
cc_918 N_A_1216_457#_M1024_g N_VPWR_c_2017_n 0.00178709f $X=7.845 $Y=2.285 $X2=0
+ $Y2=0
cc_919 N_A_1216_457#_c_1157_n N_VPWR_c_2030_n 0.0036205f $X=6.22 $Y=2.495 $X2=0
+ $Y2=0
cc_920 N_A_1216_457#_M1024_g N_VPWR_c_2010_n 9.49986e-19 $X=7.845 $Y=2.285 $X2=0
+ $Y2=0
cc_921 N_A_1216_457#_c_1157_n N_VPWR_c_2010_n 0.0045483f $X=6.22 $Y=2.495 $X2=0
+ $Y2=0
cc_922 N_A_1216_457#_c_1156_n N_A_204_119#_c_2214_n 0.0264503f $X=6.3 $Y=0.47
+ $X2=0 $Y2=0
cc_923 N_A_1216_457#_c_1156_n N_A_204_119#_c_2216_n 0.00182767f $X=6.3 $Y=0.47
+ $X2=0 $Y2=0
cc_924 N_A_1216_457#_c_1157_n N_A_204_119#_c_2216_n 0.0902162f $X=6.22 $Y=2.495
+ $X2=0 $Y2=0
cc_925 N_A_1216_457#_c_1159_n N_A_204_119#_c_2216_n 0.0129096f $X=6.3 $Y=1.11
+ $X2=0 $Y2=0
cc_926 N_A_1216_457#_c_1156_n N_A_204_119#_c_2217_n 0.0140048f $X=6.3 $Y=0.47
+ $X2=0 $Y2=0
cc_927 N_A_1216_457#_c_1156_n N_VGND_c_2459_n 0.0117747f $X=6.3 $Y=0.47 $X2=0
+ $Y2=0
cc_928 N_A_1216_457#_c_1158_n N_VGND_c_2459_n 0.0183798f $X=7.705 $Y=1.11 $X2=0
+ $Y2=0
cc_929 N_A_1216_457#_c_1156_n N_VGND_c_2470_n 0.0178561f $X=6.3 $Y=0.47 $X2=0
+ $Y2=0
cc_930 N_A_1216_457#_M1001_g N_VGND_c_2472_n 0.0035993f $X=7.815 $Y=0.555 $X2=0
+ $Y2=0
cc_931 N_A_1216_457#_M1004_d N_VGND_c_2480_n 0.0022543f $X=6.16 $Y=0.235 $X2=0
+ $Y2=0
cc_932 N_A_1216_457#_M1001_g N_VGND_c_2480_n 0.00567291f $X=7.815 $Y=0.555 $X2=0
+ $Y2=0
cc_933 N_A_1216_457#_c_1156_n N_VGND_c_2480_n 0.0124703f $X=6.3 $Y=0.47 $X2=0
+ $Y2=0
cc_934 N_A_1216_457#_M1001_g N_A_1492_47#_c_2640_n 0.00719336f $X=7.815 $Y=0.555
+ $X2=0 $Y2=0
cc_935 N_A_1216_457#_c_1158_n N_A_1492_47#_c_2640_n 0.0165877f $X=7.705 $Y=1.11
+ $X2=0 $Y2=0
cc_936 N_A_1216_457#_c_1160_n N_A_1492_47#_c_2640_n 0.00321293f $X=7.865 $Y=1.19
+ $X2=0 $Y2=0
cc_937 N_A_1216_457#_M1001_g N_A_1492_47#_c_2646_n 0.00178579f $X=7.815 $Y=0.555
+ $X2=0 $Y2=0
cc_938 N_A_1216_457#_M1001_g N_A_1492_47#_c_2639_n 0.00953562f $X=7.815 $Y=0.555
+ $X2=0 $Y2=0
cc_939 N_A_1216_457#_c_1160_n N_A_1492_47#_c_2639_n 0.0044494f $X=7.865 $Y=1.19
+ $X2=0 $Y2=0
cc_940 N_A_1650_21#_M1046_g N_A_755_106#_c_1439_n 0.00894529f $X=8.325 $Y=2.285
+ $X2=0 $Y2=0
cc_941 N_A_1650_21#_c_1257_n N_A_755_106#_M1027_g 0.00760311f $X=10.485 $Y=0.35
+ $X2=0 $Y2=0
cc_942 N_A_1650_21#_c_1259_n N_A_755_106#_M1027_g 0.00575711f $X=10.57 $Y=1
+ $X2=0 $Y2=0
cc_943 N_A_1650_21#_c_1261_n N_A_755_106#_M1027_g 0.00107279f $X=10.655 $Y=1.085
+ $X2=0 $Y2=0
cc_944 N_A_1650_21#_c_1262_n N_A_2064_453#_M1028_d 0.0105726f $X=12.5 $Y=0.915
+ $X2=-0.19 $Y2=-0.245
cc_945 N_A_1650_21#_c_1257_n N_A_2064_453#_M1009_g 0.00293582f $X=10.485 $Y=0.35
+ $X2=0 $Y2=0
cc_946 N_A_1650_21#_c_1259_n N_A_2064_453#_M1009_g 0.0130077f $X=10.57 $Y=1
+ $X2=0 $Y2=0
cc_947 N_A_1650_21#_c_1260_n N_A_2064_453#_M1009_g 0.00767481f $X=11.59 $Y=1.085
+ $X2=0 $Y2=0
cc_948 N_A_1650_21#_c_1261_n N_A_2064_453#_M1009_g 0.00342797f $X=10.655
+ $Y=1.085 $X2=0 $Y2=0
cc_949 N_A_1650_21#_c_1263_n N_A_2064_453#_M1045_g 3.45309e-19 $X=12.65 $Y=1.765
+ $X2=0 $Y2=0
cc_950 N_A_1650_21#_M1014_g N_A_2064_453#_c_1587_n 0.0154314f $X=12.32 $Y=2.675
+ $X2=0 $Y2=0
cc_951 N_A_1650_21#_c_1252_n N_A_2064_453#_c_1587_n 0.00687498f $X=12.635
+ $Y=1.785 $X2=0 $Y2=0
cc_952 N_A_1650_21#_c_1263_n N_A_2064_453#_c_1587_n 0.0185236f $X=12.65 $Y=1.765
+ $X2=0 $Y2=0
cc_953 N_A_1650_21#_c_1264_n N_A_2064_453#_c_1587_n 0.0164032f $X=12.635 $Y=1.43
+ $X2=0 $Y2=0
cc_954 N_A_1650_21#_M1000_s N_A_2064_453#_c_1602_n 0.00302884f $X=12.96 $Y=1.785
+ $X2=0 $Y2=0
cc_955 N_A_1650_21#_M1014_g N_A_2064_453#_c_1602_n 0.00986213f $X=12.32 $Y=2.675
+ $X2=0 $Y2=0
cc_956 N_A_1650_21#_c_1252_n N_A_2064_453#_c_1602_n 0.00396478f $X=12.635
+ $Y=1.785 $X2=0 $Y2=0
cc_957 N_A_1650_21#_c_1263_n N_A_2064_453#_c_1602_n 0.0385698f $X=12.65 $Y=1.765
+ $X2=0 $Y2=0
cc_958 N_A_1650_21#_c_1263_n N_A_2064_453#_c_1588_n 0.0171867f $X=12.65 $Y=1.765
+ $X2=0 $Y2=0
cc_959 N_A_1650_21#_M1014_g N_A_2064_453#_c_1638_n 0.00200231f $X=12.32 $Y=2.675
+ $X2=0 $Y2=0
cc_960 N_A_1650_21#_c_1251_n N_A_2064_453#_c_1589_n 0.00396926f $X=12.35 $Y=1
+ $X2=0 $Y2=0
cc_961 N_A_1650_21#_c_1262_n N_A_2064_453#_c_1589_n 0.0254665f $X=12.5 $Y=0.915
+ $X2=0 $Y2=0
cc_962 N_A_1650_21#_c_1264_n N_A_2064_453#_c_1589_n 0.0250585f $X=12.635 $Y=1.43
+ $X2=0 $Y2=0
cc_963 N_A_1650_21#_M1014_g N_A_2064_453#_c_1642_n 0.00519378f $X=12.32 $Y=2.675
+ $X2=0 $Y2=0
cc_964 N_A_1650_21#_c_1257_n N_A_1861_431#_M1018_d 0.00244181f $X=10.485 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_965 N_A_1650_21#_c_1251_n N_A_1861_431#_M1028_g 0.0304793f $X=12.35 $Y=1
+ $X2=0 $Y2=0
cc_966 N_A_1650_21#_c_1260_n N_A_1861_431#_M1028_g 2.64584e-19 $X=11.59 $Y=1.085
+ $X2=0 $Y2=0
cc_967 N_A_1650_21#_c_1262_n N_A_1861_431#_M1028_g 0.00857939f $X=12.5 $Y=0.915
+ $X2=0 $Y2=0
cc_968 N_A_1650_21#_c_1264_n N_A_1861_431#_M1028_g 0.00131522f $X=12.635 $Y=1.43
+ $X2=0 $Y2=0
cc_969 N_A_1650_21#_c_1266_n N_A_1861_431#_M1028_g 0.0111579f $X=11.675 $Y=0.915
+ $X2=0 $Y2=0
cc_970 N_A_1650_21#_M1014_g N_A_1861_431#_M1021_g 0.0531965f $X=12.32 $Y=2.675
+ $X2=0 $Y2=0
cc_971 N_A_1650_21#_c_1255_n N_A_1861_431#_c_1754_n 0.00734521f $X=9.445 $Y=0.86
+ $X2=0 $Y2=0
cc_972 N_A_1650_21#_c_1257_n N_A_1861_431#_c_1754_n 0.0289606f $X=10.485 $Y=0.35
+ $X2=0 $Y2=0
cc_973 N_A_1650_21#_c_1259_n N_A_1861_431#_c_1754_n 0.024269f $X=10.57 $Y=1
+ $X2=0 $Y2=0
cc_974 N_A_1650_21#_c_1259_n N_A_1861_431#_c_1755_n 0.00369987f $X=10.57 $Y=1
+ $X2=0 $Y2=0
cc_975 N_A_1650_21#_c_1261_n N_A_1861_431#_c_1755_n 0.0131397f $X=10.655
+ $Y=1.085 $X2=0 $Y2=0
cc_976 N_A_1650_21#_c_1260_n N_A_1861_431#_c_1757_n 0.0659272f $X=11.59 $Y=1.085
+ $X2=0 $Y2=0
cc_977 N_A_1650_21#_c_1261_n N_A_1861_431#_c_1757_n 0.0130771f $X=10.655
+ $Y=1.085 $X2=0 $Y2=0
cc_978 N_A_1650_21#_c_1266_n N_A_1861_431#_c_1757_n 0.0129867f $X=11.675
+ $Y=0.915 $X2=0 $Y2=0
cc_979 N_A_1650_21#_c_1252_n N_A_1861_431#_c_1760_n 2.59784e-19 $X=12.635
+ $Y=1.785 $X2=0 $Y2=0
cc_980 N_A_1650_21#_c_1252_n N_A_1861_431#_c_1761_n 0.0136143f $X=12.635
+ $Y=1.785 $X2=0 $Y2=0
cc_981 N_A_1650_21#_c_1252_n N_RESET_B_M1000_g 0.00997473f $X=12.635 $Y=1.785
+ $X2=0 $Y2=0
cc_982 N_A_1650_21#_c_1263_n N_RESET_B_M1000_g 0.00682102f $X=12.65 $Y=1.765
+ $X2=0 $Y2=0
cc_983 N_A_1650_21#_c_1264_n N_RESET_B_M1000_g 0.00138717f $X=12.635 $Y=1.43
+ $X2=0 $Y2=0
cc_984 N_A_1650_21#_c_1251_n RESET_B 0.00104562f $X=12.35 $Y=1 $X2=0 $Y2=0
cc_985 N_A_1650_21#_c_1263_n RESET_B 0.0122543f $X=12.65 $Y=1.765 $X2=0 $Y2=0
cc_986 N_A_1650_21#_c_1264_n RESET_B 0.0178558f $X=12.635 $Y=1.43 $X2=0 $Y2=0
cc_987 N_A_1650_21#_c_1268_n RESET_B 0.0137576f $X=13.105 $Y=0.815 $X2=0 $Y2=0
cc_988 N_A_1650_21#_c_1251_n N_RESET_B_c_1875_n 0.0132466f $X=12.35 $Y=1 $X2=0
+ $Y2=0
cc_989 N_A_1650_21#_c_1263_n N_RESET_B_c_1875_n 0.00126356f $X=12.65 $Y=1.765
+ $X2=0 $Y2=0
cc_990 N_A_1650_21#_c_1264_n N_RESET_B_c_1875_n 0.00160426f $X=12.635 $Y=1.43
+ $X2=0 $Y2=0
cc_991 N_A_1650_21#_c_1268_n N_RESET_B_c_1875_n 0.00115578f $X=13.105 $Y=0.815
+ $X2=0 $Y2=0
cc_992 N_A_1650_21#_c_1251_n N_RESET_B_c_1876_n 0.00227722f $X=12.35 $Y=1 $X2=0
+ $Y2=0
cc_993 N_A_1650_21#_c_1264_n N_RESET_B_c_1876_n 0.00335215f $X=12.635 $Y=1.43
+ $X2=0 $Y2=0
cc_994 N_A_1650_21#_c_1268_n N_RESET_B_c_1876_n 0.00483637f $X=13.105 $Y=0.815
+ $X2=0 $Y2=0
cc_995 N_A_1650_21#_M1046_g N_VPWR_c_2017_n 0.0119986f $X=8.325 $Y=2.285 $X2=0
+ $Y2=0
cc_996 N_A_1650_21#_M1014_g N_VPWR_c_2019_n 0.0139387f $X=12.32 $Y=2.675 $X2=0
+ $Y2=0
cc_997 N_A_1650_21#_M1014_g N_VPWR_c_2024_n 0.00486043f $X=12.32 $Y=2.675 $X2=0
+ $Y2=0
cc_998 N_A_1650_21#_M1046_g N_VPWR_c_2010_n 7.97988e-19 $X=8.325 $Y=2.285 $X2=0
+ $Y2=0
cc_999 N_A_1650_21#_M1014_g N_VPWR_c_2010_n 0.00459803f $X=12.32 $Y=2.675 $X2=0
+ $Y2=0
cc_1000 N_A_1650_21#_c_1255_n N_VGND_M1008_s 0.0031962f $X=9.445 $Y=0.86 $X2=0
+ $Y2=0
cc_1001 N_A_1650_21#_c_1248_n N_VGND_c_2460_n 0.00433715f $X=8.325 $Y=0.985
+ $X2=0 $Y2=0
cc_1002 N_A_1650_21#_c_1255_n N_VGND_c_2460_n 0.0203836f $X=9.445 $Y=0.86 $X2=0
+ $Y2=0
cc_1003 N_A_1650_21#_c_1258_n N_VGND_c_2460_n 0.00697078f $X=9.615 $Y=0.35 $X2=0
+ $Y2=0
cc_1004 N_A_1650_21#_c_1257_n N_VGND_c_2461_n 0.0128975f $X=10.485 $Y=0.35 $X2=0
+ $Y2=0
cc_1005 N_A_1650_21#_c_1259_n N_VGND_c_2461_n 0.0247537f $X=10.57 $Y=1 $X2=0
+ $Y2=0
cc_1006 N_A_1650_21#_c_1260_n N_VGND_c_2461_n 0.0259705f $X=11.59 $Y=1.085 $X2=0
+ $Y2=0
cc_1007 N_A_1650_21#_c_1268_n N_VGND_c_2462_n 0.0132651f $X=13.105 $Y=0.815
+ $X2=0 $Y2=0
cc_1008 N_A_1650_21#_c_1248_n N_VGND_c_2472_n 0.00359964f $X=8.325 $Y=0.985
+ $X2=0 $Y2=0
cc_1009 N_A_1650_21#_c_1257_n N_VGND_c_2474_n 0.06373f $X=10.485 $Y=0.35 $X2=0
+ $Y2=0
cc_1010 N_A_1650_21#_c_1258_n N_VGND_c_2474_n 0.0114622f $X=9.615 $Y=0.35 $X2=0
+ $Y2=0
cc_1011 N_A_1650_21#_c_1251_n N_VGND_c_2478_n 0.00329085f $X=12.35 $Y=1 $X2=0
+ $Y2=0
cc_1012 N_A_1650_21#_c_1268_n N_VGND_c_2478_n 0.00474015f $X=13.105 $Y=0.815
+ $X2=0 $Y2=0
cc_1013 N_A_1650_21#_c_1248_n N_VGND_c_2480_n 0.0068655f $X=8.325 $Y=0.985 $X2=0
+ $Y2=0
cc_1014 N_A_1650_21#_c_1251_n N_VGND_c_2480_n 0.00602479f $X=12.35 $Y=1 $X2=0
+ $Y2=0
cc_1015 N_A_1650_21#_c_1255_n N_VGND_c_2480_n 0.0110318f $X=9.445 $Y=0.86 $X2=0
+ $Y2=0
cc_1016 N_A_1650_21#_c_1256_n N_VGND_c_2480_n 0.00530975f $X=8.82 $Y=0.86 $X2=0
+ $Y2=0
cc_1017 N_A_1650_21#_c_1257_n N_VGND_c_2480_n 0.0383974f $X=10.485 $Y=0.35 $X2=0
+ $Y2=0
cc_1018 N_A_1650_21#_c_1258_n N_VGND_c_2480_n 0.00657784f $X=9.615 $Y=0.35 $X2=0
+ $Y2=0
cc_1019 N_A_1650_21#_c_1262_n N_VGND_c_2480_n 0.00203075f $X=12.5 $Y=0.915 $X2=0
+ $Y2=0
cc_1020 N_A_1650_21#_c_1265_n N_VGND_c_2480_n 0.00765369f $X=13.02 $Y=0.915
+ $X2=0 $Y2=0
cc_1021 N_A_1650_21#_c_1266_n N_VGND_c_2480_n 3.74539e-19 $X=11.675 $Y=0.915
+ $X2=0 $Y2=0
cc_1022 N_A_1650_21#_c_1267_n N_VGND_c_2480_n 0.00629953f $X=12.65 $Y=0.915
+ $X2=0 $Y2=0
cc_1023 N_A_1650_21#_c_1268_n N_VGND_c_2480_n 0.00729036f $X=13.105 $Y=0.815
+ $X2=0 $Y2=0
cc_1024 N_A_1650_21#_c_1256_n N_A_1492_47#_M1007_d 0.00338509f $X=8.82 $Y=0.86
+ $X2=0 $Y2=0
cc_1025 N_A_1650_21#_c_1248_n N_A_1492_47#_c_2640_n 5.86656e-19 $X=8.325
+ $Y=0.985 $X2=0 $Y2=0
cc_1026 N_A_1650_21#_c_1248_n N_A_1492_47#_c_2639_n 0.0107116f $X=8.325 $Y=0.985
+ $X2=0 $Y2=0
cc_1027 N_A_1650_21#_c_1254_n N_A_1492_47#_c_2639_n 0.00338401f $X=8.655 $Y=1.15
+ $X2=0 $Y2=0
cc_1028 N_A_1650_21#_c_1256_n N_A_1492_47#_c_2639_n 0.00829455f $X=8.82 $Y=0.86
+ $X2=0 $Y2=0
cc_1029 N_A_1650_21#_c_1255_n A_1880_57# 2.73984e-19 $X=9.445 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_1030 N_A_1650_21#_c_1406_p A_1880_57# 5.84499e-19 $X=9.53 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_1031 N_A_1650_21#_c_1258_n A_1880_57# 2.73984e-19 $X=9.615 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_1032 N_A_1650_21#_c_1259_n A_2066_101# 0.00388749f $X=10.57 $Y=1 $X2=-0.19
+ $Y2=-0.245
cc_1033 N_A_1650_21#_c_1266_n N_A_2279_57#_M1011_d 0.0014164f $X=11.675 $Y=0.915
+ $X2=-0.19 $Y2=-0.245
cc_1034 N_A_1650_21#_c_1267_n N_A_2279_57#_M1047_d 0.00262963f $X=12.65 $Y=0.915
+ $X2=0 $Y2=0
cc_1035 N_A_1650_21#_c_1251_n N_A_2279_57#_c_2669_n 0.00898335f $X=12.35 $Y=1
+ $X2=0 $Y2=0
cc_1036 N_A_1650_21#_c_1262_n N_A_2279_57#_c_2669_n 0.0169324f $X=12.5 $Y=0.915
+ $X2=0 $Y2=0
cc_1037 N_A_1650_21#_c_1266_n N_A_2279_57#_c_2669_n 0.00183465f $X=11.675
+ $Y=0.915 $X2=0 $Y2=0
cc_1038 N_A_1650_21#_c_1251_n N_A_2279_57#_c_2670_n 0.00104723f $X=12.35 $Y=1
+ $X2=0 $Y2=0
cc_1039 N_A_1650_21#_c_1260_n N_A_2279_57#_c_2670_n 0.00875866f $X=11.59
+ $Y=1.085 $X2=0 $Y2=0
cc_1040 N_A_1650_21#_c_1266_n N_A_2279_57#_c_2670_n 0.00373478f $X=11.675
+ $Y=0.915 $X2=0 $Y2=0
cc_1041 N_A_1650_21#_c_1251_n N_A_2279_57#_c_2671_n 0.00681277f $X=12.35 $Y=1
+ $X2=0 $Y2=0
cc_1042 N_A_1650_21#_c_1262_n N_A_2279_57#_c_2671_n 0.00285218f $X=12.5 $Y=0.915
+ $X2=0 $Y2=0
cc_1043 N_A_1650_21#_c_1267_n N_A_2279_57#_c_2671_n 0.0119673f $X=12.65 $Y=0.915
+ $X2=0 $Y2=0
cc_1044 N_A_1650_21#_c_1268_n N_A_2279_57#_c_2671_n 6.75592e-19 $X=13.105
+ $Y=0.815 $X2=0 $Y2=0
cc_1045 N_A_755_106#_M1027_g N_A_2064_453#_M1009_g 0.0695271f $X=10.255 $Y=0.715
+ $X2=0 $Y2=0
cc_1046 N_A_755_106#_c_1441_n N_A_2064_453#_c_1596_n 2.60863e-19 $X=10.18
+ $Y=1.77 $X2=0 $Y2=0
cc_1047 N_A_755_106#_c_1441_n N_A_2064_453#_c_1598_n 0.00625521f $X=10.18
+ $Y=1.77 $X2=0 $Y2=0
cc_1048 N_A_755_106#_M1027_g N_A_1861_431#_c_1754_n 0.0121315f $X=10.255
+ $Y=0.715 $X2=0 $Y2=0
cc_1049 N_A_755_106#_M1027_g N_A_1861_431#_c_1755_n 0.0100161f $X=10.255
+ $Y=0.715 $X2=0 $Y2=0
cc_1050 N_A_755_106#_c_1441_n N_A_1861_431#_c_1756_n 0.0071565f $X=10.18 $Y=1.77
+ $X2=0 $Y2=0
cc_1051 N_A_755_106#_M1027_g N_A_1861_431#_c_1756_n 0.00392669f $X=10.255
+ $Y=0.715 $X2=0 $Y2=0
cc_1052 N_A_755_106#_M1035_g N_A_1861_431#_c_1764_n 0.00935401f $X=9.23 $Y=2.575
+ $X2=0 $Y2=0
cc_1053 N_A_755_106#_c_1442_n N_A_1861_431#_c_1764_n 0.00402606f $X=9.54 $Y=1.77
+ $X2=0 $Y2=0
cc_1054 N_A_755_106#_c_1441_n N_A_1861_431#_c_1759_n 0.00182307f $X=10.18
+ $Y=1.77 $X2=0 $Y2=0
cc_1055 N_A_755_106#_M1027_g N_A_1861_431#_c_1759_n 0.00776443f $X=10.255
+ $Y=0.715 $X2=0 $Y2=0
cc_1056 N_A_755_106#_c_1446_n N_VPWR_c_2014_n 0.0258611f $X=4.14 $Y=2.515 $X2=0
+ $Y2=0
cc_1057 N_A_755_106#_M1042_g N_VPWR_c_2015_n 0.0148371f $X=4.915 $Y=2.605 $X2=0
+ $Y2=0
cc_1058 N_A_755_106#_c_1436_n N_VPWR_c_2015_n 0.0248025f $X=6.36 $Y=3.15 $X2=0
+ $Y2=0
cc_1059 N_A_755_106#_M1043_g N_VPWR_c_2016_n 0.00692076f $X=6.435 $Y=2.495 $X2=0
+ $Y2=0
cc_1060 N_A_755_106#_c_1439_n N_VPWR_c_2016_n 0.0252872f $X=9.155 $Y=3.15 $X2=0
+ $Y2=0
cc_1061 N_A_755_106#_c_1439_n N_VPWR_c_2017_n 0.0253854f $X=9.155 $Y=3.15 $X2=0
+ $Y2=0
cc_1062 N_A_755_106#_M1035_g N_VPWR_c_2017_n 0.00681122f $X=9.23 $Y=2.575 $X2=0
+ $Y2=0
cc_1063 N_A_755_106#_c_1437_n N_VPWR_c_2022_n 0.00763802f $X=4.99 $Y=3.15 $X2=0
+ $Y2=0
cc_1064 N_A_755_106#_c_1446_n N_VPWR_c_2022_n 0.0160569f $X=4.14 $Y=2.515 $X2=0
+ $Y2=0
cc_1065 N_A_755_106#_c_1436_n N_VPWR_c_2030_n 0.05147f $X=6.36 $Y=3.15 $X2=0
+ $Y2=0
cc_1066 N_A_755_106#_c_1439_n N_VPWR_c_2031_n 0.0348115f $X=9.155 $Y=3.15 $X2=0
+ $Y2=0
cc_1067 N_A_755_106#_c_1439_n N_VPWR_c_2032_n 0.0216899f $X=9.155 $Y=3.15 $X2=0
+ $Y2=0
cc_1068 N_A_755_106#_c_1436_n N_VPWR_c_2010_n 0.0403927f $X=6.36 $Y=3.15 $X2=0
+ $Y2=0
cc_1069 N_A_755_106#_c_1437_n N_VPWR_c_2010_n 0.01061f $X=4.99 $Y=3.15 $X2=0
+ $Y2=0
cc_1070 N_A_755_106#_c_1439_n N_VPWR_c_2010_n 0.085243f $X=9.155 $Y=3.15 $X2=0
+ $Y2=0
cc_1071 N_A_755_106#_c_1444_n N_VPWR_c_2010_n 0.00852157f $X=6.435 $Y=3.15 $X2=0
+ $Y2=0
cc_1072 N_A_755_106#_c_1446_n N_VPWR_c_2010_n 0.0109452f $X=4.14 $Y=2.515 $X2=0
+ $Y2=0
cc_1073 N_A_755_106#_c_1422_n N_A_204_119#_c_2207_n 5.9741e-19 $X=4.345 $Y=1.1
+ $X2=0 $Y2=0
cc_1074 N_A_755_106#_c_1432_n N_A_204_119#_c_2207_n 0.0145828f $X=4.05 $Y=0.79
+ $X2=0 $Y2=0
cc_1075 N_A_755_106#_c_1422_n N_A_204_119#_c_2209_n 3.36008e-19 $X=4.345 $Y=1.1
+ $X2=0 $Y2=0
cc_1076 N_A_755_106#_c_1432_n N_A_204_119#_c_2209_n 0.0284756f $X=4.05 $Y=0.79
+ $X2=0 $Y2=0
cc_1077 N_A_755_106#_c_1421_n N_A_204_119#_c_2210_n 0.00174475f $X=4.75 $Y=1.1
+ $X2=0 $Y2=0
cc_1078 N_A_755_106#_c_1422_n N_A_204_119#_c_2210_n 0.00542572f $X=4.345 $Y=1.1
+ $X2=0 $Y2=0
cc_1079 N_A_755_106#_c_1423_n N_A_204_119#_c_2210_n 0.0112231f $X=4.825 $Y=1.025
+ $X2=0 $Y2=0
cc_1080 N_A_755_106#_c_1432_n N_A_204_119#_c_2210_n 0.0281997f $X=4.05 $Y=0.79
+ $X2=0 $Y2=0
cc_1081 N_A_755_106#_c_1423_n N_A_204_119#_c_2326_n 0.0159464f $X=4.825 $Y=1.025
+ $X2=0 $Y2=0
cc_1082 N_A_755_106#_c_1428_n N_A_204_119#_c_2326_n 9.36025e-19 $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_1083 N_A_755_106#_c_1425_n N_A_204_119#_c_2212_n 0.00979455f $X=5.53 $Y=1.1
+ $X2=0 $Y2=0
cc_1084 N_A_755_106#_c_1426_n N_A_204_119#_c_2212_n 0.00747196f $X=5.605
+ $Y=1.025 $X2=0 $Y2=0
cc_1085 N_A_755_106#_c_1427_n N_A_204_119#_c_2212_n 8.34357e-19 $X=6.01 $Y=0.805
+ $X2=0 $Y2=0
cc_1086 N_A_755_106#_c_1428_n N_A_204_119#_c_2212_n 0.00474282f $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_1087 N_A_755_106#_c_1423_n N_A_204_119#_c_2213_n 0.00645431f $X=4.825
+ $Y=1.025 $X2=0 $Y2=0
cc_1088 N_A_755_106#_c_1425_n N_A_204_119#_c_2213_n 0.00130769f $X=5.53 $Y=1.1
+ $X2=0 $Y2=0
cc_1089 N_A_755_106#_c_1427_n N_A_204_119#_c_2214_n 0.0112521f $X=6.01 $Y=0.805
+ $X2=0 $Y2=0
cc_1090 N_A_755_106#_c_1429_n N_A_204_119#_c_2214_n 0.00184579f $X=6.085 $Y=0.73
+ $X2=0 $Y2=0
cc_1091 N_A_755_106#_c_1436_n N_A_204_119#_c_2221_n 0.00601418f $X=6.36 $Y=3.15
+ $X2=0 $Y2=0
cc_1092 N_A_755_106#_c_1426_n N_A_204_119#_c_2216_n 0.00534041f $X=5.605
+ $Y=1.025 $X2=0 $Y2=0
cc_1093 N_A_755_106#_c_1427_n N_A_204_119#_c_2217_n 0.00565797f $X=6.01 $Y=0.805
+ $X2=0 $Y2=0
cc_1094 N_A_755_106#_c_1423_n N_VGND_c_2458_n 0.00142601f $X=4.825 $Y=1.025
+ $X2=0 $Y2=0
cc_1095 N_A_755_106#_c_1429_n N_VGND_c_2458_n 0.00316021f $X=6.085 $Y=0.73 $X2=0
+ $Y2=0
cc_1096 N_A_755_106#_c_1423_n N_VGND_c_2468_n 7.27864e-19 $X=4.825 $Y=1.025
+ $X2=0 $Y2=0
cc_1097 N_A_755_106#_c_1427_n N_VGND_c_2470_n 0.00148975f $X=6.01 $Y=0.805 $X2=0
+ $Y2=0
cc_1098 N_A_755_106#_c_1428_n N_VGND_c_2470_n 0.0032869f $X=5.68 $Y=0.805 $X2=0
+ $Y2=0
cc_1099 N_A_755_106#_c_1429_n N_VGND_c_2470_n 0.00549284f $X=6.085 $Y=0.73 $X2=0
+ $Y2=0
cc_1100 N_A_755_106#_M1027_g N_VGND_c_2474_n 7.10185e-19 $X=10.255 $Y=0.715
+ $X2=0 $Y2=0
cc_1101 N_A_755_106#_c_1428_n N_VGND_c_2480_n 0.00555547f $X=5.68 $Y=0.805 $X2=0
+ $Y2=0
cc_1102 N_A_755_106#_c_1429_n N_VGND_c_2480_n 0.0115186f $X=6.085 $Y=0.73 $X2=0
+ $Y2=0
cc_1103 N_A_2064_453#_c_1587_n N_A_1861_431#_M1028_g 0.00153246f $X=12.235
+ $Y=2.33 $X2=0 $Y2=0
cc_1104 N_A_2064_453#_c_1589_n N_A_1861_431#_M1028_g 0.0065676f $X=12.235
+ $Y=1.37 $X2=0 $Y2=0
cc_1105 N_A_2064_453#_c_1648_p N_A_1861_431#_M1021_g 0.0091858f $X=12.15
+ $Y=2.415 $X2=0 $Y2=0
cc_1106 N_A_2064_453#_c_1587_n N_A_1861_431#_M1021_g 0.00580708f $X=12.235
+ $Y=2.33 $X2=0 $Y2=0
cc_1107 N_A_2064_453#_c_1638_n N_A_1861_431#_M1021_g 0.0111156f $X=11.685
+ $Y=2.495 $X2=0 $Y2=0
cc_1108 N_A_2064_453#_M1017_g N_A_1861_431#_c_1765_n 0.010874f $X=10.395
+ $Y=2.785 $X2=0 $Y2=0
cc_1109 N_A_2064_453#_M1009_g N_A_1861_431#_c_1754_n 3.45524e-19 $X=10.645
+ $Y=0.715 $X2=0 $Y2=0
cc_1110 N_A_2064_453#_M1009_g N_A_1861_431#_c_1755_n 0.00134715f $X=10.645
+ $Y=0.715 $X2=0 $Y2=0
cc_1111 N_A_2064_453#_M1017_g N_A_1861_431#_c_1756_n 0.00698543f $X=10.395
+ $Y=2.785 $X2=0 $Y2=0
cc_1112 N_A_2064_453#_M1009_g N_A_1861_431#_c_1756_n 0.00450783f $X=10.645
+ $Y=0.715 $X2=0 $Y2=0
cc_1113 N_A_2064_453#_c_1596_n N_A_1861_431#_c_1756_n 0.0056708f $X=10.705
+ $Y=2.265 $X2=0 $Y2=0
cc_1114 N_A_2064_453#_c_1597_n N_A_1861_431#_c_1756_n 0.0403575f $X=10.705
+ $Y=1.91 $X2=0 $Y2=0
cc_1115 N_A_2064_453#_c_1598_n N_A_1861_431#_c_1756_n 0.00697193f $X=10.705
+ $Y=1.91 $X2=0 $Y2=0
cc_1116 N_A_2064_453#_c_1600_n N_A_1861_431#_c_1756_n 0.0127199f $X=10.87
+ $Y=2.415 $X2=0 $Y2=0
cc_1117 N_A_2064_453#_M1009_g N_A_1861_431#_c_1757_n 0.011608f $X=10.645
+ $Y=0.715 $X2=0 $Y2=0
cc_1118 N_A_2064_453#_c_1597_n N_A_1861_431#_c_1757_n 0.0170708f $X=10.705
+ $Y=1.91 $X2=0 $Y2=0
cc_1119 N_A_2064_453#_c_1598_n N_A_1861_431#_c_1757_n 0.00214167f $X=10.705
+ $Y=1.91 $X2=0 $Y2=0
cc_1120 N_A_2064_453#_c_1589_n N_A_1861_431#_c_1757_n 0.0136106f $X=12.235
+ $Y=1.37 $X2=0 $Y2=0
cc_1121 N_A_2064_453#_c_1587_n N_A_1861_431#_c_1758_n 0.00692166f $X=12.235
+ $Y=2.33 $X2=0 $Y2=0
cc_1122 N_A_2064_453#_c_1589_n N_A_1861_431#_c_1758_n 9.9699e-19 $X=12.235
+ $Y=1.37 $X2=0 $Y2=0
cc_1123 N_A_2064_453#_c_1648_p N_A_1861_431#_c_1760_n 0.00564787f $X=12.15
+ $Y=2.415 $X2=0 $Y2=0
cc_1124 N_A_2064_453#_c_1587_n N_A_1861_431#_c_1760_n 0.0239776f $X=12.235
+ $Y=2.33 $X2=0 $Y2=0
cc_1125 N_A_2064_453#_c_1638_n N_A_1861_431#_c_1760_n 0.0129559f $X=11.685
+ $Y=2.495 $X2=0 $Y2=0
cc_1126 N_A_2064_453#_c_1589_n N_A_1861_431#_c_1760_n 0.00227438f $X=12.235
+ $Y=1.37 $X2=0 $Y2=0
cc_1127 N_A_2064_453#_c_1587_n N_A_1861_431#_c_1761_n 0.00349032f $X=12.235
+ $Y=2.33 $X2=0 $Y2=0
cc_1128 N_A_2064_453#_c_1638_n N_A_1861_431#_c_1761_n 0.00357324f $X=11.685
+ $Y=2.495 $X2=0 $Y2=0
cc_1129 N_A_2064_453#_c_1589_n N_A_1861_431#_c_1761_n 0.00224455f $X=12.235
+ $Y=1.37 $X2=0 $Y2=0
cc_1130 N_A_2064_453#_M1045_g N_RESET_B_M1000_g 0.0290129f $X=13.83 $Y=2.415
+ $X2=0 $Y2=0
cc_1131 N_A_2064_453#_c_1602_n N_RESET_B_M1000_g 0.0176979f $X=13.61 $Y=2.415
+ $X2=0 $Y2=0
cc_1132 N_A_2064_453#_c_1588_n N_RESET_B_M1000_g 0.0102203f $X=13.695 $Y=2.33
+ $X2=0 $Y2=0
cc_1133 N_A_2064_453#_M1036_g RESET_B 4.37111e-19 $X=13.83 $Y=0.655 $X2=0 $Y2=0
cc_1134 N_A_2064_453#_c_1590_n RESET_B 0.017367f $X=13.8 $Y=1.42 $X2=0 $Y2=0
cc_1135 N_A_2064_453#_c_1591_n RESET_B 3.13522e-19 $X=13.8 $Y=1.33 $X2=0 $Y2=0
cc_1136 N_A_2064_453#_c_1590_n N_RESET_B_c_1875_n 0.00312554f $X=13.8 $Y=1.42
+ $X2=0 $Y2=0
cc_1137 N_A_2064_453#_c_1591_n N_RESET_B_c_1875_n 0.0173645f $X=13.8 $Y=1.33
+ $X2=0 $Y2=0
cc_1138 N_A_2064_453#_M1036_g N_RESET_B_c_1876_n 0.0155103f $X=13.83 $Y=0.655
+ $X2=0 $Y2=0
cc_1139 N_A_2064_453#_M1039_g N_A_2892_137#_M1030_g 0.0150956f $X=14.82 $Y=0.895
+ $X2=0 $Y2=0
cc_1140 N_A_2064_453#_M1025_g N_A_2892_137#_M1044_g 0.0167603f $X=14.82 $Y=2.155
+ $X2=0 $Y2=0
cc_1141 N_A_2064_453#_M1036_g N_A_2892_137#_c_1910_n 0.0013742f $X=13.83
+ $Y=0.655 $X2=0 $Y2=0
cc_1142 N_A_2064_453#_c_1583_n N_A_2892_137#_c_1910_n 0.00487552f $X=14.745
+ $Y=1.33 $X2=0 $Y2=0
cc_1143 N_A_2064_453#_M1039_g N_A_2892_137#_c_1910_n 0.0114342f $X=14.82
+ $Y=0.895 $X2=0 $Y2=0
cc_1144 N_A_2064_453#_c_1586_n N_A_2892_137#_c_1910_n 9.30656e-19 $X=14.82
+ $Y=1.33 $X2=0 $Y2=0
cc_1145 N_A_2064_453#_M1045_g N_A_2892_137#_c_1915_n 0.00163362f $X=13.83
+ $Y=2.415 $X2=0 $Y2=0
cc_1146 N_A_2064_453#_M1025_g N_A_2892_137#_c_1915_n 0.0151894f $X=14.82
+ $Y=2.155 $X2=0 $Y2=0
cc_1147 N_A_2064_453#_M1025_g N_A_2892_137#_c_1911_n 0.010626f $X=14.82 $Y=2.155
+ $X2=0 $Y2=0
cc_1148 N_A_2064_453#_c_1586_n N_A_2892_137#_c_1911_n 0.00798614f $X=14.82
+ $Y=1.33 $X2=0 $Y2=0
cc_1149 N_A_2064_453#_c_1586_n N_A_2892_137#_c_1912_n 0.0213614f $X=14.82
+ $Y=1.33 $X2=0 $Y2=0
cc_1150 N_A_2064_453#_c_1583_n N_A_2892_137#_c_1913_n 0.00919862f $X=14.745
+ $Y=1.33 $X2=0 $Y2=0
cc_1151 N_A_2064_453#_M1025_g N_A_2892_137#_c_1913_n 0.00485714f $X=14.82
+ $Y=2.155 $X2=0 $Y2=0
cc_1152 N_A_2064_453#_c_1586_n N_A_2892_137#_c_1913_n 2.35411e-19 $X=14.82
+ $Y=1.33 $X2=0 $Y2=0
cc_1153 N_A_2064_453#_c_1599_n N_VPWR_M1017_d 0.00534724f $X=11.52 $Y=2.415
+ $X2=0 $Y2=0
cc_1154 N_A_2064_453#_c_1602_n N_VPWR_M1014_d 0.00645117f $X=13.61 $Y=2.415
+ $X2=0 $Y2=0
cc_1155 N_A_2064_453#_c_1602_n N_VPWR_M1000_d 0.00845321f $X=13.61 $Y=2.415
+ $X2=0 $Y2=0
cc_1156 N_A_2064_453#_c_1588_n N_VPWR_M1000_d 0.00627273f $X=13.695 $Y=2.33
+ $X2=0 $Y2=0
cc_1157 N_A_2064_453#_M1017_g N_VPWR_c_2018_n 0.00998027f $X=10.395 $Y=2.785
+ $X2=0 $Y2=0
cc_1158 N_A_2064_453#_c_1599_n N_VPWR_c_2018_n 0.0196724f $X=11.52 $Y=2.415
+ $X2=0 $Y2=0
cc_1159 N_A_2064_453#_c_1602_n N_VPWR_c_2019_n 0.0204952f $X=13.61 $Y=2.415
+ $X2=0 $Y2=0
cc_1160 N_A_2064_453#_c_1638_n N_VPWR_c_2019_n 0.0115779f $X=11.685 $Y=2.495
+ $X2=0 $Y2=0
cc_1161 N_A_2064_453#_M1045_g N_VPWR_c_2020_n 0.0104163f $X=13.83 $Y=2.415 $X2=0
+ $Y2=0
cc_1162 N_A_2064_453#_c_1602_n N_VPWR_c_2020_n 0.021264f $X=13.61 $Y=2.415 $X2=0
+ $Y2=0
cc_1163 N_A_2064_453#_M1025_g N_VPWR_c_2021_n 0.00527364f $X=14.82 $Y=2.155
+ $X2=0 $Y2=0
cc_1164 N_A_2064_453#_c_1638_n N_VPWR_c_2024_n 0.0196996f $X=11.685 $Y=2.495
+ $X2=0 $Y2=0
cc_1165 N_A_2064_453#_M1045_g N_VPWR_c_2026_n 0.00445056f $X=13.83 $Y=2.415
+ $X2=0 $Y2=0
cc_1166 N_A_2064_453#_M1025_g N_VPWR_c_2026_n 0.00312414f $X=14.82 $Y=2.155
+ $X2=0 $Y2=0
cc_1167 N_A_2064_453#_M1017_g N_VPWR_c_2032_n 0.00415733f $X=10.395 $Y=2.785
+ $X2=0 $Y2=0
cc_1168 N_A_2064_453#_M1020_d N_VPWR_c_2010_n 0.00323835f $X=11.465 $Y=2.255
+ $X2=0 $Y2=0
cc_1169 N_A_2064_453#_M1017_g N_VPWR_c_2010_n 0.00770992f $X=10.395 $Y=2.785
+ $X2=0 $Y2=0
cc_1170 N_A_2064_453#_M1045_g N_VPWR_c_2010_n 0.00899805f $X=13.83 $Y=2.415
+ $X2=0 $Y2=0
cc_1171 N_A_2064_453#_M1025_g N_VPWR_c_2010_n 0.00410284f $X=14.82 $Y=2.155
+ $X2=0 $Y2=0
cc_1172 N_A_2064_453#_c_1599_n N_VPWR_c_2010_n 0.011374f $X=11.52 $Y=2.415 $X2=0
+ $Y2=0
cc_1173 N_A_2064_453#_c_1600_n N_VPWR_c_2010_n 0.0117343f $X=10.87 $Y=2.415
+ $X2=0 $Y2=0
cc_1174 N_A_2064_453#_c_1648_p N_VPWR_c_2010_n 0.00953233f $X=12.15 $Y=2.415
+ $X2=0 $Y2=0
cc_1175 N_A_2064_453#_c_1602_n N_VPWR_c_2010_n 0.0293509f $X=13.61 $Y=2.415
+ $X2=0 $Y2=0
cc_1176 N_A_2064_453#_c_1638_n N_VPWR_c_2010_n 0.0125026f $X=11.685 $Y=2.495
+ $X2=0 $Y2=0
cc_1177 N_A_2064_453#_c_1642_n N_VPWR_c_2010_n 0.00614602f $X=12.235 $Y=2.415
+ $X2=0 $Y2=0
cc_1178 N_A_2064_453#_c_1648_p A_2395_451# 0.00679641f $X=12.15 $Y=2.415
+ $X2=-0.19 $Y2=-0.245
cc_1179 N_A_2064_453#_c_1587_n A_2395_451# 8.61155e-19 $X=12.235 $Y=2.33
+ $X2=-0.19 $Y2=-0.245
cc_1180 N_A_2064_453#_c_1642_n A_2395_451# 8.71221e-19 $X=12.235 $Y=2.415
+ $X2=-0.19 $Y2=-0.245
cc_1181 N_A_2064_453#_M1036_g N_Q_N_c_2395_n 0.00847218f $X=13.83 $Y=0.655 $X2=0
+ $Y2=0
cc_1182 N_A_2064_453#_M1039_g N_Q_N_c_2395_n 0.00366272f $X=14.82 $Y=0.895 $X2=0
+ $Y2=0
cc_1183 N_A_2064_453#_M1036_g N_Q_N_c_2396_n 0.00333139f $X=13.83 $Y=0.655 $X2=0
+ $Y2=0
cc_1184 N_A_2064_453#_c_1583_n N_Q_N_c_2396_n 0.00609999f $X=14.745 $Y=1.33
+ $X2=0 $Y2=0
cc_1185 N_A_2064_453#_c_1590_n N_Q_N_c_2396_n 0.00407834f $X=13.8 $Y=1.42 $X2=0
+ $Y2=0
cc_1186 N_A_2064_453#_M1045_g N_Q_N_c_2398_n 0.00453744f $X=13.83 $Y=2.415 $X2=0
+ $Y2=0
cc_1187 N_A_2064_453#_c_1583_n N_Q_N_c_2398_n 0.00620508f $X=14.745 $Y=1.33
+ $X2=0 $Y2=0
cc_1188 N_A_2064_453#_c_1588_n N_Q_N_c_2398_n 0.0190254f $X=13.695 $Y=2.33 $X2=0
+ $Y2=0
cc_1189 N_A_2064_453#_M1036_g N_Q_N_c_2397_n 0.00411273f $X=13.83 $Y=0.655 $X2=0
+ $Y2=0
cc_1190 N_A_2064_453#_M1045_g N_Q_N_c_2397_n 0.00251684f $X=13.83 $Y=2.415 $X2=0
+ $Y2=0
cc_1191 N_A_2064_453#_c_1583_n N_Q_N_c_2397_n 0.0148071f $X=14.745 $Y=1.33 $X2=0
+ $Y2=0
cc_1192 N_A_2064_453#_M1025_g N_Q_N_c_2397_n 0.00318595f $X=14.82 $Y=2.155 $X2=0
+ $Y2=0
cc_1193 N_A_2064_453#_c_1588_n N_Q_N_c_2397_n 0.00524694f $X=13.695 $Y=2.33
+ $X2=0 $Y2=0
cc_1194 N_A_2064_453#_c_1590_n N_Q_N_c_2397_n 0.0232923f $X=13.8 $Y=1.42 $X2=0
+ $Y2=0
cc_1195 N_A_2064_453#_c_1591_n N_Q_N_c_2397_n 0.00124625f $X=13.8 $Y=1.33 $X2=0
+ $Y2=0
cc_1196 N_A_2064_453#_M1025_g Q_N 0.00197803f $X=14.82 $Y=2.155 $X2=0 $Y2=0
cc_1197 N_A_2064_453#_M1009_g N_VGND_c_2461_n 0.00412411f $X=10.645 $Y=0.715
+ $X2=0 $Y2=0
cc_1198 N_A_2064_453#_M1036_g N_VGND_c_2462_n 0.00483983f $X=13.83 $Y=0.655
+ $X2=0 $Y2=0
cc_1199 N_A_2064_453#_c_1590_n N_VGND_c_2462_n 0.0054544f $X=13.8 $Y=1.42 $X2=0
+ $Y2=0
cc_1200 N_A_2064_453#_c_1591_n N_VGND_c_2462_n 0.00141917f $X=13.8 $Y=1.33 $X2=0
+ $Y2=0
cc_1201 N_A_2064_453#_M1039_g N_VGND_c_2463_n 0.00412273f $X=14.82 $Y=0.895
+ $X2=0 $Y2=0
cc_1202 N_A_2064_453#_M1009_g N_VGND_c_2474_n 0.00250138f $X=10.645 $Y=0.715
+ $X2=0 $Y2=0
cc_1203 N_A_2064_453#_M1036_g N_VGND_c_2476_n 0.00549284f $X=13.83 $Y=0.655
+ $X2=0 $Y2=0
cc_1204 N_A_2064_453#_M1039_g N_VGND_c_2476_n 0.00371502f $X=14.82 $Y=0.895
+ $X2=0 $Y2=0
cc_1205 N_A_2064_453#_M1009_g N_VGND_c_2480_n 0.0021835f $X=10.645 $Y=0.715
+ $X2=0 $Y2=0
cc_1206 N_A_2064_453#_M1036_g N_VGND_c_2480_n 0.0123926f $X=13.83 $Y=0.655 $X2=0
+ $Y2=0
cc_1207 N_A_2064_453#_M1039_g N_VGND_c_2480_n 0.00453162f $X=14.82 $Y=0.895
+ $X2=0 $Y2=0
cc_1208 N_A_2064_453#_M1028_d N_A_2279_57#_c_2669_n 0.00609737f $X=11.825
+ $Y=0.285 $X2=0 $Y2=0
cc_1209 N_A_1861_431#_c_1764_n N_VPWR_c_2017_n 0.012279f $X=9.445 $Y=2.68 $X2=0
+ $Y2=0
cc_1210 N_A_1861_431#_M1021_g N_VPWR_c_2018_n 0.00110178f $X=11.9 $Y=2.675 $X2=0
+ $Y2=0
cc_1211 N_A_1861_431#_c_1765_n N_VPWR_c_2018_n 0.00253202f $X=10.225 $Y=2.68
+ $X2=0 $Y2=0
cc_1212 N_A_1861_431#_M1021_g N_VPWR_c_2019_n 0.00231553f $X=11.9 $Y=2.675 $X2=0
+ $Y2=0
cc_1213 N_A_1861_431#_M1021_g N_VPWR_c_2024_n 0.00549284f $X=11.9 $Y=2.675 $X2=0
+ $Y2=0
cc_1214 N_A_1861_431#_c_1765_n N_VPWR_c_2032_n 0.0145628f $X=10.225 $Y=2.68
+ $X2=0 $Y2=0
cc_1215 N_A_1861_431#_c_1764_n N_VPWR_c_2032_n 0.0163606f $X=9.445 $Y=2.68 $X2=0
+ $Y2=0
cc_1216 N_A_1861_431#_M1021_g N_VPWR_c_2010_n 0.00645497f $X=11.9 $Y=2.675 $X2=0
+ $Y2=0
cc_1217 N_A_1861_431#_c_1765_n N_VPWR_c_2010_n 0.0228284f $X=10.225 $Y=2.68
+ $X2=0 $Y2=0
cc_1218 N_A_1861_431#_c_1764_n N_VPWR_c_2010_n 0.0120693f $X=9.445 $Y=2.68 $X2=0
+ $Y2=0
cc_1219 N_A_1861_431#_c_1765_n A_1963_515# 0.0118326f $X=10.225 $Y=2.68
+ $X2=-0.19 $Y2=-0.245
cc_1220 N_A_1861_431#_c_1756_n A_1963_515# 2.69964e-19 $X=10.31 $Y=2.595
+ $X2=-0.19 $Y2=-0.245
cc_1221 N_A_1861_431#_M1028_g N_VGND_c_2478_n 0.00329085f $X=11.75 $Y=0.605
+ $X2=0 $Y2=0
cc_1222 N_A_1861_431#_M1028_g N_VGND_c_2480_n 0.00513344f $X=11.75 $Y=0.605
+ $X2=0 $Y2=0
cc_1223 N_A_1861_431#_M1028_g N_A_2279_57#_c_2669_n 0.00892812f $X=11.75
+ $Y=0.605 $X2=0 $Y2=0
cc_1224 N_A_1861_431#_M1028_g N_A_2279_57#_c_2670_n 0.00612536f $X=11.75
+ $Y=0.605 $X2=0 $Y2=0
cc_1225 N_A_1861_431#_M1028_g N_A_2279_57#_c_2671_n 0.00105028f $X=11.75
+ $Y=0.605 $X2=0 $Y2=0
cc_1226 N_RESET_B_M1000_g N_VPWR_c_2033_n 0.00294244f $X=13.32 $Y=2.105 $X2=0
+ $Y2=0
cc_1227 N_RESET_B_M1000_g N_VPWR_c_2010_n 0.00398527f $X=13.32 $Y=2.105 $X2=0
+ $Y2=0
cc_1228 N_RESET_B_c_1876_n N_Q_N_c_2395_n 4.65727e-19 $X=13.23 $Y=1.185 $X2=0
+ $Y2=0
cc_1229 N_RESET_B_c_1876_n N_VGND_c_2462_n 0.00490885f $X=13.23 $Y=1.185 $X2=0
+ $Y2=0
cc_1230 N_RESET_B_c_1876_n N_VGND_c_2478_n 0.00385415f $X=13.23 $Y=1.185 $X2=0
+ $Y2=0
cc_1231 N_RESET_B_c_1876_n N_VGND_c_2480_n 0.0046122f $X=13.23 $Y=1.185 $X2=0
+ $Y2=0
cc_1232 N_RESET_B_c_1876_n N_A_2279_57#_c_2671_n 0.00259994f $X=13.23 $Y=1.185
+ $X2=0 $Y2=0
cc_1233 N_A_2892_137#_M1044_g N_VPWR_c_2021_n 0.00698192f $X=15.33 $Y=2.465
+ $X2=0 $Y2=0
cc_1234 N_A_2892_137#_c_1915_n N_VPWR_c_2021_n 0.0248129f $X=14.605 $Y=1.98
+ $X2=0 $Y2=0
cc_1235 N_A_2892_137#_c_1911_n N_VPWR_c_2021_n 0.0206753f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1236 N_A_2892_137#_c_1912_n N_VPWR_c_2021_n 0.002179f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1237 N_A_2892_137#_M1044_g N_VPWR_c_2034_n 0.00549284f $X=15.33 $Y=2.465
+ $X2=0 $Y2=0
cc_1238 N_A_2892_137#_M1044_g N_VPWR_c_2010_n 0.012057f $X=15.33 $Y=2.465 $X2=0
+ $Y2=0
cc_1239 N_A_2892_137#_c_1915_n N_VPWR_c_2010_n 0.00972751f $X=14.605 $Y=1.98
+ $X2=0 $Y2=0
cc_1240 N_A_2892_137#_c_1910_n N_Q_N_c_2395_n 0.0448528f $X=14.605 $Y=0.895
+ $X2=0 $Y2=0
cc_1241 N_A_2892_137#_c_1915_n N_Q_N_c_2397_n 0.0606527f $X=14.605 $Y=1.98 $X2=0
+ $Y2=0
cc_1242 N_A_2892_137#_c_1913_n N_Q_N_c_2397_n 0.0235744f $X=14.645 $Y=1.47 $X2=0
+ $Y2=0
cc_1243 N_A_2892_137#_M1044_g N_Q_c_2432_n 0.0144708f $X=15.33 $Y=2.465 $X2=0
+ $Y2=0
cc_1244 N_A_2892_137#_M1044_g N_Q_c_2433_n 0.00287652f $X=15.33 $Y=2.465 $X2=0
+ $Y2=0
cc_1245 N_A_2892_137#_c_1911_n N_Q_c_2433_n 0.00144832f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1246 N_A_2892_137#_c_1912_n N_Q_c_2433_n 0.00131892f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1247 N_A_2892_137#_M1030_g N_Q_c_2429_n 0.00440999f $X=15.33 $Y=0.685 $X2=0
+ $Y2=0
cc_1248 N_A_2892_137#_M1044_g N_Q_c_2429_n 0.00440999f $X=15.33 $Y=2.465 $X2=0
+ $Y2=0
cc_1249 N_A_2892_137#_c_1911_n N_Q_c_2429_n 0.0250957f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1250 N_A_2892_137#_c_1912_n N_Q_c_2429_n 0.00768695f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1251 N_A_2892_137#_M1030_g Q 0.00287652f $X=15.33 $Y=0.685 $X2=0 $Y2=0
cc_1252 N_A_2892_137#_c_1911_n Q 0.00144832f $X=15.27 $Y=1.47 $X2=0 $Y2=0
cc_1253 N_A_2892_137#_c_1912_n Q 0.00131892f $X=15.27 $Y=1.47 $X2=0 $Y2=0
cc_1254 N_A_2892_137#_M1030_g N_Q_c_2431_n 0.010297f $X=15.33 $Y=0.685 $X2=0
+ $Y2=0
cc_1255 N_A_2892_137#_M1030_g N_VGND_c_2463_n 0.0055345f $X=15.33 $Y=0.685 $X2=0
+ $Y2=0
cc_1256 N_A_2892_137#_c_1910_n N_VGND_c_2463_n 0.0172562f $X=14.605 $Y=0.895
+ $X2=0 $Y2=0
cc_1257 N_A_2892_137#_c_1911_n N_VGND_c_2463_n 0.0206753f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1258 N_A_2892_137#_c_1912_n N_VGND_c_2463_n 0.002179f $X=15.27 $Y=1.47 $X2=0
+ $Y2=0
cc_1259 N_A_2892_137#_c_1910_n N_VGND_c_2476_n 0.00467036f $X=14.605 $Y=0.895
+ $X2=0 $Y2=0
cc_1260 N_A_2892_137#_M1030_g N_VGND_c_2479_n 0.00520813f $X=15.33 $Y=0.685
+ $X2=0 $Y2=0
cc_1261 N_A_2892_137#_M1030_g N_VGND_c_2480_n 0.0115561f $X=15.33 $Y=0.685 $X2=0
+ $Y2=0
cc_1262 N_A_2892_137#_c_1910_n N_VGND_c_2480_n 0.00733137f $X=14.605 $Y=0.895
+ $X2=0 $Y2=0
cc_1263 N_A_27_481#_c_1960_n N_VPWR_c_2011_n 0.0240561f $X=0.28 $Y=2.55 $X2=0
+ $Y2=0
cc_1264 N_A_27_481#_c_1961_n N_VPWR_c_2011_n 0.0241543f $X=1.135 $Y=2.15 $X2=0
+ $Y2=0
cc_1265 N_A_27_481#_c_1965_n N_VPWR_c_2011_n 0.00161266f $X=1.305 $Y=2.98 $X2=0
+ $Y2=0
cc_1266 N_A_27_481#_c_1964_n N_VPWR_c_2012_n 0.0119251f $X=1.995 $Y=2.98 $X2=0
+ $Y2=0
cc_1267 N_A_27_481#_c_1966_n N_VPWR_c_2012_n 0.0336423f $X=2.16 $Y=2.55 $X2=0
+ $Y2=0
cc_1268 N_A_27_481#_c_1960_n N_VPWR_c_2028_n 0.0220321f $X=0.28 $Y=2.55 $X2=0
+ $Y2=0
cc_1269 N_A_27_481#_c_1964_n N_VPWR_c_2029_n 0.063174f $X=1.995 $Y=2.98 $X2=0
+ $Y2=0
cc_1270 N_A_27_481#_c_1965_n N_VPWR_c_2029_n 0.0114622f $X=1.305 $Y=2.98 $X2=0
+ $Y2=0
cc_1271 N_A_27_481#_c_1960_n N_VPWR_c_2010_n 0.0125808f $X=0.28 $Y=2.55 $X2=0
+ $Y2=0
cc_1272 N_A_27_481#_c_1964_n N_VPWR_c_2010_n 0.0371744f $X=1.995 $Y=2.98 $X2=0
+ $Y2=0
cc_1273 N_A_27_481#_c_1965_n N_VPWR_c_2010_n 0.00657784f $X=1.305 $Y=2.98 $X2=0
+ $Y2=0
cc_1274 N_A_27_481#_c_1963_n A_224_481# 0.00213724f $X=1.22 $Y=2.895 $X2=-0.19
+ $Y2=1.655
cc_1275 N_A_27_481#_c_1964_n N_A_204_119#_M1005_d 0.00180746f $X=1.995 $Y=2.98
+ $X2=0 $Y2=0
cc_1276 N_A_27_481#_c_1961_n N_A_204_119#_c_2218_n 0.00242297f $X=1.135 $Y=2.15
+ $X2=0 $Y2=0
cc_1277 N_A_27_481#_c_1963_n N_A_204_119#_c_2218_n 0.0232745f $X=1.22 $Y=2.895
+ $X2=0 $Y2=0
cc_1278 N_A_27_481#_c_1964_n N_A_204_119#_c_2218_n 0.0149073f $X=1.995 $Y=2.98
+ $X2=0 $Y2=0
cc_1279 N_A_27_481#_c_1966_n N_A_204_119#_c_2218_n 0.0125869f $X=2.16 $Y=2.55
+ $X2=0 $Y2=0
cc_1280 N_A_27_481#_c_1961_n N_A_204_119#_c_2220_n 0.0118379f $X=1.135 $Y=2.15
+ $X2=0 $Y2=0
cc_1281 N_A_27_481#_c_1966_n N_A_204_119#_c_2220_n 0.0115162f $X=2.16 $Y=2.55
+ $X2=0 $Y2=0
cc_1282 N_VPWR_c_2015_n N_A_204_119#_c_2221_n 0.029279f $X=5.21 $Y=2.43 $X2=0
+ $Y2=0
cc_1283 N_VPWR_c_2030_n N_A_204_119#_c_2221_n 0.00691124f $X=6.955 $Y=3.33 $X2=0
+ $Y2=0
cc_1284 N_VPWR_c_2010_n N_A_204_119#_c_2221_n 0.0087658f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1285 N_VPWR_c_2010_n A_2395_451# 0.00392033f $X=15.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1286 N_VPWR_c_2020_n Q_N 0.0145666f $X=13.615 $Y=2.87 $X2=0 $Y2=0
cc_1287 N_VPWR_c_2021_n Q_N 0.0186234f $X=15.115 $Y=1.98 $X2=0 $Y2=0
cc_1288 N_VPWR_c_2026_n Q_N 0.0238008f $X=14.95 $Y=3.33 $X2=0 $Y2=0
cc_1289 N_VPWR_c_2010_n Q_N 0.0136587f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1290 N_VPWR_c_2010_n N_Q_M1044_d 0.0023218f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1291 N_VPWR_c_2034_n N_Q_c_2432_n 0.022455f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1292 N_VPWR_c_2010_n N_Q_c_2432_n 0.0140558f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1293 N_VPWR_c_2021_n N_Q_c_2433_n 0.0462846f $X=15.115 $Y=1.98 $X2=0 $Y2=0
cc_1294 N_A_204_119#_c_2203_n N_VGND_M1003_d 0.00403103f $X=2.3 $Y=1.175 $X2=0
+ $Y2=0
cc_1295 N_A_204_119#_c_2210_n N_VGND_M1022_d 0.00107963f $X=4.875 $Y=0.35 $X2=0
+ $Y2=0
cc_1296 N_A_204_119#_c_2326_n N_VGND_M1022_d 0.00552863f $X=4.96 $Y=0.83 $X2=0
+ $Y2=0
cc_1297 N_A_204_119#_c_2212_n N_VGND_M1022_d 0.0074493f $X=5.705 $Y=0.915 $X2=0
+ $Y2=0
cc_1298 N_A_204_119#_c_2199_n N_VGND_c_2455_n 0.0145731f $X=1.16 $Y=0.805 $X2=0
+ $Y2=0
cc_1299 N_A_204_119#_c_2199_n N_VGND_c_2456_n 0.0137594f $X=1.16 $Y=0.805 $X2=0
+ $Y2=0
cc_1300 N_A_204_119#_c_2200_n N_VGND_c_2456_n 0.016113f $X=1.975 $Y=1.26 $X2=0
+ $Y2=0
cc_1301 N_A_204_119#_c_2203_n N_VGND_c_2456_n 0.0405564f $X=2.3 $Y=1.175 $X2=0
+ $Y2=0
cc_1302 N_A_204_119#_c_2205_n N_VGND_c_2456_n 0.0141592f $X=2.385 $Y=0.35 $X2=0
+ $Y2=0
cc_1303 N_A_204_119#_c_2204_n N_VGND_c_2457_n 0.0137879f $X=2.915 $Y=0.35 $X2=0
+ $Y2=0
cc_1304 N_A_204_119#_c_2206_n N_VGND_c_2457_n 0.0380885f $X=3 $Y=1.15 $X2=0
+ $Y2=0
cc_1305 N_A_204_119#_c_2207_n N_VGND_c_2457_n 0.0136257f $X=3.615 $Y=1.235 $X2=0
+ $Y2=0
cc_1306 N_A_204_119#_c_2209_n N_VGND_c_2457_n 0.0228252f $X=3.7 $Y=1.15 $X2=0
+ $Y2=0
cc_1307 N_A_204_119#_c_2211_n N_VGND_c_2457_n 0.0137873f $X=3.785 $Y=0.35 $X2=0
+ $Y2=0
cc_1308 N_A_204_119#_c_2210_n N_VGND_c_2458_n 0.0138501f $X=4.875 $Y=0.35 $X2=0
+ $Y2=0
cc_1309 N_A_204_119#_c_2326_n N_VGND_c_2458_n 0.0153766f $X=4.96 $Y=0.83 $X2=0
+ $Y2=0
cc_1310 N_A_204_119#_c_2212_n N_VGND_c_2458_n 0.0182058f $X=5.705 $Y=0.915 $X2=0
+ $Y2=0
cc_1311 N_A_204_119#_c_2214_n N_VGND_c_2458_n 0.024888f $X=5.87 $Y=0.47 $X2=0
+ $Y2=0
cc_1312 N_A_204_119#_c_2199_n N_VGND_c_2464_n 0.0074415f $X=1.16 $Y=0.805 $X2=0
+ $Y2=0
cc_1313 N_A_204_119#_c_2204_n N_VGND_c_2466_n 0.0431887f $X=2.915 $Y=0.35 $X2=0
+ $Y2=0
cc_1314 N_A_204_119#_c_2205_n N_VGND_c_2466_n 0.011374f $X=2.385 $Y=0.35 $X2=0
+ $Y2=0
cc_1315 N_A_204_119#_c_2210_n N_VGND_c_2468_n 0.0774992f $X=4.875 $Y=0.35 $X2=0
+ $Y2=0
cc_1316 N_A_204_119#_c_2211_n N_VGND_c_2468_n 0.0114622f $X=3.785 $Y=0.35 $X2=0
+ $Y2=0
cc_1317 N_A_204_119#_c_2214_n N_VGND_c_2470_n 0.0163773f $X=5.87 $Y=0.47 $X2=0
+ $Y2=0
cc_1318 N_A_204_119#_M1004_s N_VGND_c_2480_n 0.00297283f $X=5.725 $Y=0.235 $X2=0
+ $Y2=0
cc_1319 N_A_204_119#_c_2199_n N_VGND_c_2480_n 0.00902447f $X=1.16 $Y=0.805 $X2=0
+ $Y2=0
cc_1320 N_A_204_119#_c_2204_n N_VGND_c_2480_n 0.0258056f $X=2.915 $Y=0.35 $X2=0
+ $Y2=0
cc_1321 N_A_204_119#_c_2205_n N_VGND_c_2480_n 0.00585508f $X=2.385 $Y=0.35 $X2=0
+ $Y2=0
cc_1322 N_A_204_119#_c_2210_n N_VGND_c_2480_n 0.0473062f $X=4.875 $Y=0.35 $X2=0
+ $Y2=0
cc_1323 N_A_204_119#_c_2211_n N_VGND_c_2480_n 0.00657784f $X=3.785 $Y=0.35 $X2=0
+ $Y2=0
cc_1324 N_A_204_119#_c_2212_n N_VGND_c_2480_n 0.0145562f $X=5.705 $Y=0.915 $X2=0
+ $Y2=0
cc_1325 N_A_204_119#_c_2214_n N_VGND_c_2480_n 0.00959046f $X=5.87 $Y=0.47 $X2=0
+ $Y2=0
cc_1326 N_Q_N_c_2395_n N_VGND_c_2463_n 0.0132665f $X=14.045 $Y=0.43 $X2=0 $Y2=0
cc_1327 N_Q_N_c_2395_n N_VGND_c_2476_n 0.0268376f $X=14.045 $Y=0.43 $X2=0 $Y2=0
cc_1328 N_Q_N_M1036_d N_VGND_c_2480_n 0.0023218f $X=13.905 $Y=0.235 $X2=0 $Y2=0
cc_1329 N_Q_N_c_2395_n N_VGND_c_2480_n 0.0165708f $X=14.045 $Y=0.43 $X2=0 $Y2=0
cc_1330 N_Q_c_2431_n N_VGND_c_2463_n 0.0320595f $X=15.545 $Y=0.43 $X2=0 $Y2=0
cc_1331 N_Q_c_2431_n N_VGND_c_2479_n 0.022455f $X=15.545 $Y=0.43 $X2=0 $Y2=0
cc_1332 N_Q_c_2431_n N_VGND_c_2480_n 0.0141183f $X=15.545 $Y=0.43 $X2=0 $Y2=0
cc_1333 N_VGND_c_2480_n A_1318_47# 0.00899413f $X=15.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1334 N_VGND_c_2480_n N_A_1492_47#_M1026_d 0.0022543f $X=15.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1335 N_VGND_c_2480_n N_A_1492_47#_M1007_d 0.00232217f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1336 N_VGND_c_2472_n N_A_1492_47#_c_2646_n 0.017823f $X=8.935 $Y=0 $X2=0
+ $Y2=0
cc_1337 N_VGND_c_2480_n N_A_1492_47#_c_2646_n 0.0124841f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1338 N_VGND_c_2460_n N_A_1492_47#_c_2639_n 0.0141648f $X=9.1 $Y=0.47 $X2=0
+ $Y2=0
cc_1339 N_VGND_c_2472_n N_A_1492_47#_c_2639_n 0.0514925f $X=8.935 $Y=0 $X2=0
+ $Y2=0
cc_1340 N_VGND_c_2480_n N_A_1492_47#_c_2639_n 0.0339233f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1341 N_VGND_c_2478_n N_A_2279_57#_c_2669_n 0.0417281f $X=13.45 $Y=0 $X2=0
+ $Y2=0
cc_1342 N_VGND_c_2480_n N_A_2279_57#_c_2669_n 0.0250167f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1343 N_VGND_c_2461_n N_A_2279_57#_c_2670_n 0.0145581f $X=11.025 $Y=0.54 $X2=0
+ $Y2=0
cc_1344 N_VGND_c_2478_n N_A_2279_57#_c_2670_n 0.0210491f $X=13.45 $Y=0 $X2=0
+ $Y2=0
cc_1345 N_VGND_c_2480_n N_A_2279_57#_c_2670_n 0.0122835f $X=15.6 $Y=0 $X2=0
+ $Y2=0
cc_1346 N_VGND_c_2478_n N_A_2279_57#_c_2671_n 0.0159546f $X=13.45 $Y=0 $X2=0
+ $Y2=0
cc_1347 N_VGND_c_2480_n N_A_2279_57#_c_2671_n 0.00934402f $X=15.6 $Y=0 $X2=0
+ $Y2=0
