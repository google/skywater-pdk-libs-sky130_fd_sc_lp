* NGSPICE file created from sky130_fd_sc_lp__and4_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4_1 A B C D VGND VNB VPB VPWR X
M1000 VGND D a_327_47# VNB nshort w=420000u l=150000u
+  ad=2.835e+11p pd=2.46e+06u as=1.638e+11p ps=1.62e+06u
M1001 a_123_47# A a_40_47# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.113e+11p ps=1.37e+06u
M1002 a_219_47# B a_123_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1003 VPWR B a_40_47# VPB phighvt w=420000u l=150000u
+  ad=7.854e+11p pd=6.88e+06u as=2.814e+11p ps=3.02e+06u
M1004 VPWR D a_40_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_40_47# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1006 a_327_47# C a_219_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_40_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1008 a_40_47# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_40_47# C VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

