* File: sky130_fd_sc_lp__fa_4.pxi.spice
* Created: Fri Aug 28 10:35:00 2020
* 
x_PM_SKY130_FD_SC_LP__FA_4%A N_A_c_190_n N_A_M1038_g N_A_M1030_g N_A_M1016_g
+ N_A_M1006_g N_A_M1035_g N_A_M1031_g N_A_M1003_g N_A_M1029_g N_A_c_211_n
+ N_A_c_196_n N_A_c_197_n N_A_c_213_n N_A_c_214_n N_A_c_215_n N_A_c_216_n
+ N_A_c_217_n N_A_c_198_n N_A_c_219_n N_A_c_220_n N_A_c_199_n N_A_c_200_n
+ N_A_c_201_n N_A_c_202_n N_A_c_203_n N_A_c_204_n N_A_c_205_n A A A
+ PM_SKY130_FD_SC_LP__FA_4%A
x_PM_SKY130_FD_SC_LP__FA_4%A_328_131# N_A_328_131#_M1025_d N_A_328_131#_M1024_d
+ N_A_328_131#_M1039_g N_A_328_131#_M1012_g N_A_328_131#_c_395_n
+ N_A_328_131#_M1014_g N_A_328_131#_M1010_g N_A_328_131#_c_397_n
+ N_A_328_131#_M1015_g N_A_328_131#_M1022_g N_A_328_131#_c_399_n
+ N_A_328_131#_M1034_g N_A_328_131#_M1023_g N_A_328_131#_c_401_n
+ N_A_328_131#_M1036_g N_A_328_131#_M1037_g N_A_328_131#_c_427_n
+ N_A_328_131#_c_420_n N_A_328_131#_c_429_n N_A_328_131#_c_403_n
+ N_A_328_131#_c_404_n N_A_328_131#_c_405_n N_A_328_131#_c_406_n
+ N_A_328_131#_c_407_n N_A_328_131#_c_408_n N_A_328_131#_c_409_n
+ N_A_328_131#_c_410_n N_A_328_131#_c_411_n N_A_328_131#_c_412_n
+ N_A_328_131#_c_413_n N_A_328_131#_c_414_n PM_SKY130_FD_SC_LP__FA_4%A_328_131#
x_PM_SKY130_FD_SC_LP__FA_4%CIN N_CIN_M1025_g N_CIN_M1024_g N_CIN_c_598_n
+ N_CIN_M1032_g N_CIN_M1026_g N_CIN_c_600_n N_CIN_M1001_g N_CIN_M1007_g
+ N_CIN_c_602_n CIN CIN CIN N_CIN_c_604_n PM_SKY130_FD_SC_LP__FA_4%CIN
x_PM_SKY130_FD_SC_LP__FA_4%B N_B_M1011_g N_B_M1005_g N_B_c_696_n N_B_c_697_n
+ N_B_M1028_g N_B_M1019_g N_B_c_700_n N_B_M1033_g N_B_M1009_g N_B_c_702_n
+ N_B_M1008_g N_B_M1002_g N_B_c_704_n N_B_c_705_n N_B_c_706_n B B N_B_c_694_n
+ PM_SKY130_FD_SC_LP__FA_4%B
x_PM_SKY130_FD_SC_LP__FA_4%A_884_131# N_A_884_131#_M1039_d N_A_884_131#_M1012_d
+ N_A_884_131#_M1004_g N_A_884_131#_M1000_g N_A_884_131#_M1017_g
+ N_A_884_131#_M1013_g N_A_884_131#_M1018_g N_A_884_131#_M1020_g
+ N_A_884_131#_M1021_g N_A_884_131#_M1027_g N_A_884_131#_c_842_n
+ N_A_884_131#_c_846_n N_A_884_131#_c_830_n N_A_884_131#_c_831_n
+ N_A_884_131#_c_872_n N_A_884_131#_c_839_n N_A_884_131#_c_832_n
+ N_A_884_131#_c_833_n PM_SKY130_FD_SC_LP__FA_4%A_884_131#
x_PM_SKY130_FD_SC_LP__FA_4%A_27_440# N_A_27_440#_M1038_s N_A_27_440#_M1011_d
+ N_A_27_440#_c_956_n N_A_27_440#_c_957_n N_A_27_440#_c_963_n
+ N_A_27_440#_c_966_n PM_SKY130_FD_SC_LP__FA_4%A_27_440#
x_PM_SKY130_FD_SC_LP__FA_4%VPWR N_VPWR_M1038_d N_VPWR_M1006_d N_VPWR_M1009_d
+ N_VPWR_M1029_d N_VPWR_M1013_d N_VPWR_M1027_d N_VPWR_M1022_d N_VPWR_M1037_d
+ N_VPWR_c_981_n N_VPWR_c_982_n N_VPWR_c_983_n N_VPWR_c_984_n N_VPWR_c_985_n
+ N_VPWR_c_986_n N_VPWR_c_987_n N_VPWR_c_988_n N_VPWR_c_989_n N_VPWR_c_990_n
+ N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_993_n N_VPWR_c_994_n N_VPWR_c_995_n
+ VPWR N_VPWR_c_996_n N_VPWR_c_997_n N_VPWR_c_998_n N_VPWR_c_999_n
+ N_VPWR_c_1000_n N_VPWR_c_1001_n N_VPWR_c_1002_n N_VPWR_c_1003_n
+ N_VPWR_c_1004_n N_VPWR_c_980_n PM_SKY130_FD_SC_LP__FA_4%VPWR
x_PM_SKY130_FD_SC_LP__FA_4%A_604_419# N_A_604_419#_M1026_d N_A_604_419#_M1031_d
+ N_A_604_419#_c_1124_n N_A_604_419#_c_1122_n N_A_604_419#_c_1123_n
+ PM_SKY130_FD_SC_LP__FA_4%A_604_419#
x_PM_SKY130_FD_SC_LP__FA_4%SUM N_SUM_M1004_d N_SUM_M1018_d N_SUM_M1000_s
+ N_SUM_M1020_s N_SUM_c_1207_p N_SUM_c_1194_n N_SUM_c_1149_n N_SUM_c_1150_n
+ N_SUM_c_1153_n N_SUM_c_1154_n N_SUM_c_1208_p N_SUM_c_1198_n N_SUM_c_1151_n SUM
+ SUM PM_SKY130_FD_SC_LP__FA_4%SUM
x_PM_SKY130_FD_SC_LP__FA_4%COUT N_COUT_M1014_s N_COUT_M1034_s N_COUT_M1010_s
+ N_COUT_M1023_s N_COUT_c_1263_p N_COUT_c_1247_n N_COUT_c_1220_n N_COUT_c_1224_n
+ N_COUT_c_1215_n N_COUT_c_1216_n N_COUT_c_1264_p N_COUT_c_1251_n
+ N_COUT_c_1235_n N_COUT_c_1217_n N_COUT_c_1239_n N_COUT_c_1218_n COUT COUT COUT
+ PM_SKY130_FD_SC_LP__FA_4%COUT
x_PM_SKY130_FD_SC_LP__FA_4%A_37_131# N_A_37_131#_M1030_s N_A_37_131#_M1005_d
+ N_A_37_131#_c_1295_p N_A_37_131#_c_1272_n N_A_37_131#_c_1273_n
+ N_A_37_131#_c_1274_n PM_SKY130_FD_SC_LP__FA_4%A_37_131#
x_PM_SKY130_FD_SC_LP__FA_4%VGND N_VGND_M1030_d N_VGND_M1016_d N_VGND_M1033_d
+ N_VGND_M1003_d N_VGND_M1017_s N_VGND_M1021_s N_VGND_M1015_d N_VGND_M1036_d
+ N_VGND_c_1297_n N_VGND_c_1298_n N_VGND_c_1299_n N_VGND_c_1300_n
+ N_VGND_c_1301_n N_VGND_c_1302_n N_VGND_c_1303_n N_VGND_c_1304_n
+ N_VGND_c_1305_n N_VGND_c_1306_n N_VGND_c_1307_n N_VGND_c_1308_n
+ N_VGND_c_1309_n N_VGND_c_1310_n N_VGND_c_1311_n VGND N_VGND_c_1312_n
+ N_VGND_c_1313_n N_VGND_c_1314_n N_VGND_c_1315_n N_VGND_c_1316_n
+ N_VGND_c_1317_n N_VGND_c_1318_n N_VGND_c_1319_n N_VGND_c_1320_n
+ N_VGND_c_1321_n PM_SKY130_FD_SC_LP__FA_4%VGND
x_PM_SKY130_FD_SC_LP__FA_4%A_604_131# N_A_604_131#_M1032_d N_A_604_131#_M1035_d
+ N_A_604_131#_c_1449_n N_A_604_131#_c_1435_n N_A_604_131#_c_1436_n
+ N_A_604_131#_c_1451_n PM_SKY130_FD_SC_LP__FA_4%A_604_131#
cc_1 VNB N_A_c_190_n 0.011219f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.87
cc_2 VNB N_A_M1030_g 0.0360524f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.865
cc_3 VNB N_A_M1016_g 0.0195724f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.865
cc_4 VNB N_A_M1006_g 0.00271254f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=2.415
cc_5 VNB N_A_M1035_g 0.0344149f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=0.865
cc_6 VNB N_A_M1003_g 0.025938f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=0.865
cc_7 VNB N_A_c_196_n 0.00315819f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.535
cc_8 VNB N_A_c_197_n 0.0224752f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.535
cc_9 VNB N_A_c_198_n 8.21569e-19 $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=1.915
cc_10 VNB N_A_c_199_n 0.00114733f $X=-0.19 $Y=-0.245 $X2=4.995 $Y2=1.51
cc_11 VNB N_A_c_200_n 0.00234961f $X=-0.19 $Y=-0.245 $X2=5.625 $Y2=1.51
cc_12 VNB N_A_c_201_n 0.0255557f $X=-0.19 $Y=-0.245 $X2=5.625 $Y2=1.51
cc_13 VNB N_A_c_202_n 0.031869f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.43
cc_14 VNB N_A_c_203_n 0.00688227f $X=-0.19 $Y=-0.245 $X2=3.725 $Y2=1.65
cc_15 VNB N_A_c_204_n 0.00791757f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.77
cc_16 VNB N_A_c_205_n 0.0030075f $X=-0.19 $Y=-0.245 $X2=3.99 $Y2=1.65
cc_17 VNB N_A_328_131#_M1039_g 0.0220843f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.865
cc_18 VNB N_A_328_131#_M1012_g 4.99233e-19 $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.865
cc_19 VNB N_A_328_131#_c_395_n 0.0160639f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.595
cc_20 VNB N_A_328_131#_M1010_g 0.00726984f $X=-0.19 $Y=-0.245 $X2=3.915
+ $Y2=0.865
cc_21 VNB N_A_328_131#_c_397_n 0.0158822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_328_131#_M1022_g 0.00706662f $X=-0.19 $Y=-0.245 $X2=5.535
+ $Y2=1.345
cc_23 VNB N_A_328_131#_c_399_n 0.0158799f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=0.865
cc_24 VNB N_A_328_131#_M1023_g 0.00706364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_328_131#_c_401_n 0.0183577f $X=-0.19 $Y=-0.245 $X2=0.477 $Y2=1.93
cc_26 VNB N_A_328_131#_M1037_g 0.00760894f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=2.015
cc_27 VNB N_A_328_131#_c_403_n 0.0012359f $X=-0.19 $Y=-0.245 $X2=5.625 $Y2=1.51
cc_28 VNB N_A_328_131#_c_404_n 0.0293644f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.65
cc_29 VNB N_A_328_131#_c_405_n 0.00170639f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.43
cc_30 VNB N_A_328_131#_c_406_n 0.0286244f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.43
cc_31 VNB N_A_328_131#_c_407_n 0.00312262f $X=-0.19 $Y=-0.245 $X2=3.725 $Y2=1.65
cc_32 VNB N_A_328_131#_c_408_n 0.020465f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.65
cc_33 VNB N_A_328_131#_c_409_n 0.00570196f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.77
cc_34 VNB N_A_328_131#_c_410_n 0.00464823f $X=-0.19 $Y=-0.245 $X2=4.91 $Y2=1.51
cc_35 VNB N_A_328_131#_c_411_n 0.00632307f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_36 VNB N_A_328_131#_c_412_n 0.0025015f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.58
cc_37 VNB N_A_328_131#_c_413_n 0.00909559f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.65
cc_38 VNB N_A_328_131#_c_414_n 0.080058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_CIN_M1025_g 0.0365703f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.04
cc_40 VNB N_CIN_c_598_n 0.0831098f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.37
cc_41 VNB N_CIN_M1032_g 0.050607f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.265
cc_42 VNB N_CIN_c_600_n 0.140163f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.595
cc_43 VNB N_CIN_M1001_g 0.0590722f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=1.605
cc_44 VNB N_CIN_c_602_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=1.935
cc_45 VNB CIN 0.0185594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_CIN_c_604_n 0.0477663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_B_M1005_g 0.0356388f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.37
cc_48 VNB N_B_M1028_g 0.0326938f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.865
cc_49 VNB N_B_M1033_g 0.0365621f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=1.935
cc_50 VNB N_B_M1008_g 0.0341419f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.675
cc_51 VNB B 0.00674178f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.015
cc_52 VNB N_B_c_694_n 0.0173544f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=2.985
cc_53 VNB N_A_884_131#_M1004_g 0.0243689f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.865
cc_54 VNB N_A_884_131#_M1000_g 4.07161e-19 $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.865
cc_55 VNB N_A_884_131#_M1017_g 0.0205741f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=2.415
cc_56 VNB N_A_884_131#_M1013_g 4.56879e-19 $X=-0.19 $Y=-0.245 $X2=3.915
+ $Y2=0.865
cc_57 VNB N_A_884_131#_M1018_g 0.0205741f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=2.415
cc_58 VNB N_A_884_131#_M1020_g 4.55536e-19 $X=-0.19 $Y=-0.245 $X2=5.535
+ $Y2=0.865
cc_59 VNB N_A_884_131#_M1021_g 0.0205233f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=2.415
cc_60 VNB N_A_884_131#_M1027_g 3.83102e-19 $X=-0.19 $Y=-0.245 $X2=0.477
+ $Y2=1.535
cc_61 VNB N_A_884_131#_c_830_n 0.00334161f $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=2.895
cc_62 VNB N_A_884_131#_c_831_n 5.19797e-19 $X=-0.19 $Y=-0.245 $X2=3.99 $Y2=1.83
cc_63 VNB N_A_884_131#_c_832_n 0.00101481f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.65
cc_64 VNB N_A_884_131#_c_833_n 0.0758761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VPWR_c_980_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_SUM_c_1149_n 0.00244912f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=1.935
cc_67 VNB N_SUM_c_1150_n 0.00176422f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=2.415
cc_68 VNB N_SUM_c_1151_n 0.00240549f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.535
cc_69 VNB SUM 0.003435f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.535
cc_70 VNB COUT 0.00781009f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.895
cc_71 VNB COUT 0.0318513f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=2.985
cc_72 VNB N_A_37_131#_c_1272_n 0.00692019f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=1.265
cc_73 VNB N_A_37_131#_c_1273_n 0.00987073f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.865
cc_74 VNB N_A_37_131#_c_1274_n 0.00485103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1297_n 0.0219084f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.345
cc_76 VNB N_VGND_c_1298_n 0.00827229f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.675
cc_77 VNB N_VGND_c_1299_n 0.0156201f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=2.04
cc_78 VNB N_VGND_c_1300_n 0.0142618f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.535
cc_79 VNB N_VGND_c_1301_n 3.12649e-19 $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.1
cc_80 VNB N_VGND_c_1302_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=1.915
cc_81 VNB N_VGND_c_1303_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=4.995 $Y2=1.51
cc_82 VNB N_VGND_c_1304_n 0.0105251f $X=-0.19 $Y=-0.245 $X2=5.625 $Y2=1.51
cc_83 VNB N_VGND_c_1305_n 0.0197167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1306_n 0.0559241f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.43
cc_85 VNB N_VGND_c_1307_n 0.00522339f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.43
cc_86 VNB N_VGND_c_1308_n 0.0135019f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.65
cc_87 VNB N_VGND_c_1309_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.77
cc_88 VNB N_VGND_c_1310_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=3.99 $Y2=1.65
cc_89 VNB N_VGND_c_1311_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=4.91 $Y2=1.51
cc_90 VNB N_VGND_c_1312_n 0.0196742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1313_n 0.0366836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1314_n 0.020195f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.605
cc_93 VNB N_VGND_c_1315_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1316_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1317_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1318_n 0.00476075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1319_n 0.00476075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1320_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1321_n 0.474157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_604_131#_c_1435_n 0.00681158f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=1.265
cc_101 VNB N_A_604_131#_c_1436_n 0.00330771f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.865
cc_102 VPB N_A_c_190_n 0.0210602f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=1.87
cc_103 VPB N_A_M1038_g 0.0260509f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.52
cc_104 VPB N_A_M1006_g 0.0278277f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=2.415
cc_105 VPB N_A_M1031_g 0.0190357f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=2.415
cc_106 VPB N_A_M1029_g 0.0352262f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=2.415
cc_107 VPB N_A_c_211_n 0.0199875f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=2.04
cc_108 VPB N_A_c_196_n 0.00244919f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.535
cc_109 VPB N_A_c_213_n 0.0136976f $X=-0.19 $Y=1.655 $X2=1.5 $Y2=2.015
cc_110 VPB N_A_c_214_n 0.0046376f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.015
cc_111 VPB N_A_c_215_n 0.00192254f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.895
cc_112 VPB N_A_c_216_n 0.0153529f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.985
cc_113 VPB N_A_c_217_n 0.00283663f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=2.985
cc_114 VPB N_A_c_198_n 0.00163811f $X=-0.19 $Y=1.655 $X2=2.38 $Y2=1.915
cc_115 VPB N_A_c_219_n 0.00264829f $X=-0.19 $Y=1.655 $X2=2.38 $Y2=2.895
cc_116 VPB N_A_c_220_n 0.0118117f $X=-0.19 $Y=1.655 $X2=4.825 $Y2=1.83
cc_117 VPB N_A_c_199_n 0.00325724f $X=-0.19 $Y=1.655 $X2=4.995 $Y2=1.51
cc_118 VPB N_A_c_200_n 0.00428754f $X=-0.19 $Y=1.655 $X2=5.625 $Y2=1.51
cc_119 VPB N_A_c_201_n 0.00645089f $X=-0.19 $Y=1.655 $X2=5.625 $Y2=1.51
cc_120 VPB N_A_c_203_n 0.00958993f $X=-0.19 $Y=1.655 $X2=3.725 $Y2=1.65
cc_121 VPB N_A_c_204_n 0.0209832f $X=-0.19 $Y=1.655 $X2=3.825 $Y2=1.77
cc_122 VPB N_A_c_205_n 0.00111665f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=1.65
cc_123 VPB N_A_328_131#_M1012_g 0.0323198f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.865
cc_124 VPB N_A_328_131#_M1010_g 0.0198609f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=0.865
cc_125 VPB N_A_328_131#_M1022_g 0.0189123f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.345
cc_126 VPB N_A_328_131#_M1023_g 0.0188927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_328_131#_M1037_g 0.0224628f $X=-0.19 $Y=1.655 $X2=1.5 $Y2=2.015
cc_128 VPB N_A_328_131#_c_420_n 0.00146803f $X=-0.19 $Y=1.655 $X2=2.38 $Y2=1.915
cc_129 VPB N_A_328_131#_c_405_n 0.00134016f $X=-0.19 $Y=1.655 $X2=2.445 $Y2=1.43
cc_130 VPB N_CIN_M1025_g 0.0353446f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.04
cc_131 VPB N_CIN_M1032_g 0.0304888f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=1.265
cc_132 VPB N_CIN_M1001_g 0.0299283f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=1.605
cc_133 VPB N_B_M1011_g 0.0304658f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.52
cc_134 VPB N_B_c_696_n 0.0783488f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.865
cc_135 VPB N_B_c_697_n 0.011606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_B_M1028_g 0.00912762f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.865
cc_137 VPB N_B_M1019_g 0.0236363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_B_c_700_n 0.0745387f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=1.605
cc_139 VPB N_B_M1033_g 0.0414402f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=1.935
cc_140 VPB N_B_c_702_n 0.130142f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.345
cc_141 VPB N_B_M1008_g 0.0463653f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.675
cc_142 VPB N_B_c_704_n 0.0221681f $X=-0.19 $Y=1.655 $X2=0.477 $Y2=1.535
cc_143 VPB N_B_c_705_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.535
cc_144 VPB N_B_c_706_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB B 0.00722357f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.015
cc_146 VPB N_B_c_694_n 0.0183533f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=2.985
cc_147 VPB N_A_884_131#_M1000_g 0.0215558f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.865
cc_148 VPB N_A_884_131#_M1013_g 0.0187403f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=0.865
cc_149 VPB N_A_884_131#_M1020_g 0.0187396f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=0.865
cc_150 VPB N_A_884_131#_M1027_g 0.0180652f $X=-0.19 $Y=1.655 $X2=0.477 $Y2=1.535
cc_151 VPB N_A_884_131#_c_831_n 0.00178693f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=1.83
cc_152 VPB N_A_884_131#_c_839_n 0.00462762f $X=-0.19 $Y=1.655 $X2=3.725 $Y2=1.65
cc_153 VPB N_A_27_440#_c_956_n 0.0183797f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.37
cc_154 VPB N_A_27_440#_c_957_n 0.0177123f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.865
cc_155 VPB N_VPWR_c_981_n 0.00700827f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.345
cc_156 VPB N_VPWR_c_982_n 0.00696865f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.675
cc_157 VPB N_VPWR_c_983_n 0.0140274f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=2.04
cc_158 VPB N_VPWR_c_984_n 0.00772441f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.535
cc_159 VPB N_VPWR_c_985_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.985
cc_160 VPB N_VPWR_c_986_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=4.995 $Y2=1.51
cc_161 VPB N_VPWR_c_987_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=2.412 $Y2=1.59
cc_162 VPB N_VPWR_c_988_n 0.0104993f $X=-0.19 $Y=1.655 $X2=3.825 $Y2=1.65
cc_163 VPB N_VPWR_c_989_n 0.0412086f $X=-0.19 $Y=1.655 $X2=3.825 $Y2=1.77
cc_164 VPB N_VPWR_c_990_n 0.0569084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_991_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.58
cc_166 VPB N_VPWR_c_992_n 0.0129398f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.58
cc_167 VPB N_VPWR_c_993_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_994_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_995_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=1.535
cc_170 VPB N_VPWR_c_996_n 0.0173493f $X=-0.19 $Y=1.655 $X2=2.445 $Y2=1.265
cc_171 VPB N_VPWR_c_997_n 0.0444797f $X=-0.19 $Y=1.655 $X2=5.625 $Y2=1.51
cc_172 VPB N_VPWR_c_998_n 0.016463f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=1.65
cc_173 VPB N_VPWR_c_999_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1000_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1001_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1002_n 0.00290382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1003_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1004_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_980_n 0.0674705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_604_419#_c_1122_n 0.00444837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_604_419#_c_1123_n 0.00397285f $X=-0.19 $Y=1.655 $X2=2.51
+ $Y2=2.415
cc_182 VPB N_SUM_c_1153_n 0.00282821f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=2.415
cc_183 VPB N_SUM_c_1154_n 0.00202208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB SUM 0.00305599f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.535
cc_185 VPB N_COUT_c_1215_n 0.00348586f $X=-0.19 $Y=1.655 $X2=3.915 $Y2=2.415
cc_186 VPB N_COUT_c_1216_n 0.00232154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_COUT_c_1217_n 0.0110982f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.535
cc_188 VPB N_COUT_c_1218_n 0.00167091f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.015
cc_189 VPB COUT 0.00499244f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.985
cc_190 N_A_M1035_g N_A_328_131#_M1039_g 0.0201657f $X=3.915 $Y=0.865 $X2=0 $Y2=0
cc_191 N_A_c_220_n N_A_328_131#_M1012_g 0.0151795f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_192 N_A_c_199_n N_A_328_131#_M1012_g 6.09211e-19 $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_193 N_A_c_204_n N_A_328_131#_M1012_g 0.0268146f $X=3.825 $Y=1.77 $X2=0 $Y2=0
cc_194 N_A_c_205_n N_A_328_131#_M1012_g 6.18426e-19 $X=3.99 $Y=1.65 $X2=0 $Y2=0
cc_195 N_A_M1016_g N_A_328_131#_c_427_n 0.00148156f $X=2.355 $Y=0.865 $X2=0
+ $Y2=0
cc_196 N_A_c_213_n N_A_328_131#_c_420_n 0.00364168f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_197 N_A_c_216_n N_A_328_131#_c_429_n 0.018719f $X=2.295 $Y=2.985 $X2=0 $Y2=0
cc_198 N_A_M1035_g N_A_328_131#_c_403_n 2.40744e-19 $X=3.915 $Y=0.865 $X2=0
+ $Y2=0
cc_199 N_A_c_220_n N_A_328_131#_c_403_n 0.0181821f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_200 N_A_c_205_n N_A_328_131#_c_403_n 0.0124292f $X=3.99 $Y=1.65 $X2=0 $Y2=0
cc_201 N_A_M1035_g N_A_328_131#_c_404_n 0.0214835f $X=3.915 $Y=0.865 $X2=0 $Y2=0
cc_202 N_A_c_220_n N_A_328_131#_c_404_n 0.0043992f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_203 N_A_c_199_n N_A_328_131#_c_404_n 6.21665e-19 $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_204 N_A_c_205_n N_A_328_131#_c_404_n 7.30355e-19 $X=3.99 $Y=1.65 $X2=0 $Y2=0
cc_205 N_A_M1006_g N_A_328_131#_c_405_n 0.00132453f $X=2.51 $Y=2.415 $X2=0 $Y2=0
cc_206 N_A_c_213_n N_A_328_131#_c_405_n 0.00431188f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_207 N_A_c_219_n N_A_328_131#_c_405_n 0.0565547f $X=2.38 $Y=2.895 $X2=0 $Y2=0
cc_208 N_A_c_202_n N_A_328_131#_c_405_n 0.00141615f $X=2.445 $Y=1.43 $X2=0 $Y2=0
cc_209 N_A_M1016_g N_A_328_131#_c_406_n 0.00653813f $X=2.355 $Y=0.865 $X2=0
+ $Y2=0
cc_210 N_A_M1035_g N_A_328_131#_c_406_n 0.00532943f $X=3.915 $Y=0.865 $X2=0
+ $Y2=0
cc_211 N_A_c_198_n N_A_328_131#_c_406_n 0.020835f $X=2.38 $Y=1.915 $X2=0 $Y2=0
cc_212 N_A_c_220_n N_A_328_131#_c_406_n 0.00534362f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_213 N_A_c_202_n N_A_328_131#_c_406_n 0.00380655f $X=2.445 $Y=1.43 $X2=0 $Y2=0
cc_214 N_A_c_203_n N_A_328_131#_c_406_n 0.0519393f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_215 N_A_c_198_n N_A_328_131#_c_407_n 6.92306e-19 $X=2.38 $Y=1.915 $X2=0 $Y2=0
cc_216 N_A_M1003_g N_A_328_131#_c_408_n 0.00313943f $X=5.535 $Y=0.865 $X2=0
+ $Y2=0
cc_217 N_A_c_220_n N_A_328_131#_c_408_n 0.00381913f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_218 N_A_c_199_n N_A_328_131#_c_408_n 0.0104605f $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_219 N_A_c_200_n N_A_328_131#_c_408_n 0.0425097f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_220 N_A_c_201_n N_A_328_131#_c_408_n 0.00449089f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_221 N_A_c_220_n N_A_328_131#_c_409_n 0.00328682f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_222 N_A_c_199_n N_A_328_131#_c_409_n 0.00133914f $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_223 N_A_M1016_g N_A_328_131#_c_410_n 0.00141615f $X=2.355 $Y=0.865 $X2=0
+ $Y2=0
cc_224 N_A_c_198_n N_A_328_131#_c_410_n 0.0499916f $X=2.38 $Y=1.915 $X2=0 $Y2=0
cc_225 N_A_M1035_g N_A_328_131#_c_411_n 4.41668e-19 $X=3.915 $Y=0.865 $X2=0
+ $Y2=0
cc_226 N_A_c_220_n N_A_328_131#_c_411_n 0.0132745f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_227 N_A_c_199_n N_A_328_131#_c_411_n 0.0160106f $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_c_213_n N_CIN_M1025_g 0.00959991f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_229 N_A_c_215_n N_CIN_M1025_g 0.0249334f $X=1.585 $Y=2.895 $X2=0 $Y2=0
cc_230 N_A_M1016_g N_CIN_c_598_n 0.00910836f $X=2.355 $Y=0.865 $X2=0 $Y2=0
cc_231 N_A_M1016_g N_CIN_M1032_g 0.012712f $X=2.355 $Y=0.865 $X2=0 $Y2=0
cc_232 N_A_M1006_g N_CIN_M1032_g 0.0265433f $X=2.51 $Y=2.415 $X2=0 $Y2=0
cc_233 N_A_c_198_n N_CIN_M1032_g 9.53603e-19 $X=2.38 $Y=1.915 $X2=0 $Y2=0
cc_234 N_A_c_219_n N_CIN_M1032_g 0.00111652f $X=2.38 $Y=2.895 $X2=0 $Y2=0
cc_235 N_A_c_202_n N_CIN_M1032_g 0.0169959f $X=2.445 $Y=1.43 $X2=0 $Y2=0
cc_236 N_A_c_203_n N_CIN_M1032_g 0.0296894f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_237 N_A_M1035_g N_CIN_c_600_n 0.00912852f $X=3.915 $Y=0.865 $X2=0 $Y2=0
cc_238 N_A_c_220_n N_CIN_M1001_g 0.00688654f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_239 N_A_c_199_n N_CIN_M1001_g 0.0121476f $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_240 N_A_c_200_n N_CIN_M1001_g 3.52512e-19 $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_241 N_A_M1016_g CIN 8.7152e-19 $X=2.355 $Y=0.865 $X2=0 $Y2=0
cc_242 N_A_c_190_n N_B_M1011_g 0.0152587f $X=0.43 $Y=1.87 $X2=0 $Y2=0
cc_243 N_A_M1038_g N_B_M1011_g 0.0278636f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_244 N_A_c_213_n N_B_M1011_g 0.0125405f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_245 N_A_c_215_n N_B_M1011_g 0.00241398f $X=1.585 $Y=2.895 $X2=0 $Y2=0
cc_246 N_A_c_217_n N_B_M1011_g 0.00153144f $X=1.67 $Y=2.985 $X2=0 $Y2=0
cc_247 N_A_M1030_g N_B_M1005_g 0.0258248f $X=0.525 $Y=0.865 $X2=0 $Y2=0
cc_248 N_A_c_196_n N_B_M1005_g 0.00217389f $X=0.425 $Y=1.535 $X2=0 $Y2=0
cc_249 N_A_c_216_n N_B_c_696_n 0.0074072f $X=2.295 $Y=2.985 $X2=0 $Y2=0
cc_250 N_A_c_217_n N_B_c_696_n 0.00186329f $X=1.67 $Y=2.985 $X2=0 $Y2=0
cc_251 N_A_M1016_g N_B_M1028_g 0.0652132f $X=2.355 $Y=0.865 $X2=0 $Y2=0
cc_252 N_A_M1006_g N_B_M1028_g 0.00755688f $X=2.51 $Y=2.415 $X2=0 $Y2=0
cc_253 N_A_c_198_n N_B_M1028_g 0.00136049f $X=2.38 $Y=1.915 $X2=0 $Y2=0
cc_254 N_A_c_215_n N_B_M1019_g 0.00151717f $X=1.585 $Y=2.895 $X2=0 $Y2=0
cc_255 N_A_c_216_n N_B_M1019_g 0.0147428f $X=2.295 $Y=2.985 $X2=0 $Y2=0
cc_256 N_A_M1006_g N_B_c_700_n 0.0102834f $X=2.51 $Y=2.415 $X2=0 $Y2=0
cc_257 N_A_c_216_n N_B_c_700_n 0.00461574f $X=2.295 $Y=2.985 $X2=0 $Y2=0
cc_258 N_A_M1035_g N_B_M1033_g 0.0262059f $X=3.915 $Y=0.865 $X2=0 $Y2=0
cc_259 N_A_M1031_g N_B_M1033_g 0.0164487f $X=3.915 $Y=2.415 $X2=0 $Y2=0
cc_260 N_A_c_203_n N_B_M1033_g 0.0238282f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_261 N_A_c_204_n N_B_M1033_g 0.0214417f $X=3.825 $Y=1.77 $X2=0 $Y2=0
cc_262 N_A_M1031_g N_B_c_702_n 0.0103719f $X=3.915 $Y=2.415 $X2=0 $Y2=0
cc_263 N_A_M1003_g N_B_M1008_g 0.149922f $X=5.535 $Y=0.865 $X2=0 $Y2=0
cc_264 N_A_c_199_n N_B_M1008_g 0.00553966f $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_265 N_A_c_200_n N_B_M1008_g 0.0144842f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_266 N_A_M1006_g N_B_c_704_n 0.0610771f $X=2.51 $Y=2.415 $X2=0 $Y2=0
cc_267 N_A_c_213_n N_B_c_704_n 4.17085e-19 $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_268 N_A_c_198_n N_B_c_704_n 6.18804e-19 $X=2.38 $Y=1.915 $X2=0 $Y2=0
cc_269 N_A_c_219_n N_B_c_704_n 0.00739179f $X=2.38 $Y=2.895 $X2=0 $Y2=0
cc_270 N_A_c_196_n B 0.0166584f $X=0.425 $Y=1.535 $X2=0 $Y2=0
cc_271 N_A_c_213_n B 0.0576538f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_272 N_A_c_196_n N_B_c_694_n 0.00730401f $X=0.425 $Y=1.535 $X2=0 $Y2=0
cc_273 N_A_c_197_n N_B_c_694_n 0.0152587f $X=0.425 $Y=1.535 $X2=0 $Y2=0
cc_274 N_A_c_213_n N_B_c_694_n 0.00604771f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_275 N_A_M1003_g N_A_884_131#_M1004_g 0.0199525f $X=5.535 $Y=0.865 $X2=0 $Y2=0
cc_276 N_A_M1029_g N_A_884_131#_M1000_g 0.0218227f $X=5.535 $Y=2.415 $X2=0 $Y2=0
cc_277 N_A_M1003_g N_A_884_131#_c_842_n 0.0185022f $X=5.535 $Y=0.865 $X2=0 $Y2=0
cc_278 N_A_c_199_n N_A_884_131#_c_842_n 0.00472841f $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_279 N_A_c_200_n N_A_884_131#_c_842_n 0.0199051f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_280 N_A_c_201_n N_A_884_131#_c_842_n 0.00345804f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_281 N_A_M1029_g N_A_884_131#_c_846_n 0.0162967f $X=5.535 $Y=2.415 $X2=0 $Y2=0
cc_282 N_A_c_220_n N_A_884_131#_c_846_n 0.00514713f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_283 N_A_c_199_n N_A_884_131#_c_846_n 0.0107671f $X=4.995 $Y=1.51 $X2=0 $Y2=0
cc_284 N_A_c_200_n N_A_884_131#_c_846_n 0.023006f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_285 N_A_c_201_n N_A_884_131#_c_846_n 0.00389275f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_286 N_A_M1003_g N_A_884_131#_c_830_n 0.00544585f $X=5.535 $Y=0.865 $X2=0
+ $Y2=0
cc_287 N_A_c_200_n N_A_884_131#_c_830_n 0.00366138f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_288 N_A_c_201_n N_A_884_131#_c_830_n 3.12813e-19 $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_289 N_A_M1029_g N_A_884_131#_c_831_n 0.00809794f $X=5.535 $Y=2.415 $X2=0
+ $Y2=0
cc_290 N_A_c_200_n N_A_884_131#_c_831_n 0.0086723f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_291 N_A_c_201_n N_A_884_131#_c_831_n 7.38926e-19 $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_292 N_A_c_220_n N_A_884_131#_c_839_n 0.0204173f $X=4.825 $Y=1.83 $X2=0 $Y2=0
cc_293 N_A_c_200_n N_A_884_131#_c_832_n 0.0151549f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_294 N_A_c_201_n N_A_884_131#_c_832_n 0.00128858f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_295 N_A_c_200_n N_A_884_131#_c_833_n 2.96928e-19 $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_296 N_A_c_201_n N_A_884_131#_c_833_n 0.0169107f $X=5.625 $Y=1.51 $X2=0 $Y2=0
cc_297 N_A_c_213_n N_A_27_440#_M1011_d 0.00686599f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_298 N_A_M1038_g N_A_27_440#_c_956_n 8.05401e-19 $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_299 N_A_c_211_n N_A_27_440#_c_956_n 0.00263051f $X=0.43 $Y=2.04 $X2=0 $Y2=0
cc_300 N_A_c_214_n N_A_27_440#_c_956_n 0.00828741f $X=0.695 $Y=2.015 $X2=0 $Y2=0
cc_301 N_A_M1038_g N_A_27_440#_c_957_n 2.20346e-19 $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_302 N_A_M1038_g N_A_27_440#_c_963_n 0.0123659f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_303 N_A_c_213_n N_A_27_440#_c_963_n 0.0244873f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_304 N_A_c_214_n N_A_27_440#_c_963_n 0.0191347f $X=0.695 $Y=2.015 $X2=0 $Y2=0
cc_305 N_A_c_213_n N_A_27_440#_c_966_n 0.0153048f $X=1.5 $Y=2.015 $X2=0 $Y2=0
cc_306 N_A_c_215_n N_A_27_440#_c_966_n 0.0225376f $X=1.585 $Y=2.895 $X2=0 $Y2=0
cc_307 N_A_M1038_g N_VPWR_c_981_n 0.0100889f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_308 N_A_c_215_n N_VPWR_c_981_n 0.00656286f $X=1.585 $Y=2.895 $X2=0 $Y2=0
cc_309 N_A_c_217_n N_VPWR_c_981_n 0.00551624f $X=1.67 $Y=2.985 $X2=0 $Y2=0
cc_310 N_A_M1006_g N_VPWR_c_982_n 9.45943e-19 $X=2.51 $Y=2.415 $X2=0 $Y2=0
cc_311 N_A_c_216_n N_VPWR_c_982_n 0.0154744f $X=2.295 $Y=2.985 $X2=0 $Y2=0
cc_312 N_A_c_219_n N_VPWR_c_982_n 0.0330704f $X=2.38 $Y=2.895 $X2=0 $Y2=0
cc_313 N_A_c_203_n N_VPWR_c_982_n 0.0161129f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_314 N_A_M1031_g N_VPWR_c_983_n 0.00321833f $X=3.915 $Y=2.415 $X2=0 $Y2=0
cc_315 N_A_M1029_g N_VPWR_c_984_n 0.0114426f $X=5.535 $Y=2.415 $X2=0 $Y2=0
cc_316 N_A_M1029_g N_VPWR_c_990_n 0.00431487f $X=5.535 $Y=2.415 $X2=0 $Y2=0
cc_317 N_A_M1038_g N_VPWR_c_996_n 0.00410575f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_318 N_A_c_216_n N_VPWR_c_997_n 0.0515041f $X=2.295 $Y=2.985 $X2=0 $Y2=0
cc_319 N_A_c_217_n N_VPWR_c_997_n 0.0115893f $X=1.67 $Y=2.985 $X2=0 $Y2=0
cc_320 N_A_M1038_g N_VPWR_c_980_n 0.00427039f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_321 N_A_M1006_g N_VPWR_c_980_n 7.53851e-19 $X=2.51 $Y=2.415 $X2=0 $Y2=0
cc_322 N_A_M1031_g N_VPWR_c_980_n 9.39239e-19 $X=3.915 $Y=2.415 $X2=0 $Y2=0
cc_323 N_A_M1029_g N_VPWR_c_980_n 0.00477801f $X=5.535 $Y=2.415 $X2=0 $Y2=0
cc_324 N_A_c_216_n N_VPWR_c_980_n 0.0267156f $X=2.295 $Y=2.985 $X2=0 $Y2=0
cc_325 N_A_c_217_n N_VPWR_c_980_n 0.00583135f $X=1.67 $Y=2.985 $X2=0 $Y2=0
cc_326 N_A_c_219_n A_445_419# 0.00538035f $X=2.38 $Y=2.895 $X2=-0.19 $Y2=-0.245
cc_327 N_A_M1031_g N_A_604_419#_c_1124_n 0.0125876f $X=3.915 $Y=2.415 $X2=0
+ $Y2=0
cc_328 N_A_c_203_n N_A_604_419#_c_1124_n 0.0470971f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_329 N_A_c_204_n N_A_604_419#_c_1124_n 0.00397056f $X=3.825 $Y=1.77 $X2=0
+ $Y2=0
cc_330 N_A_c_203_n N_A_604_419#_c_1122_n 0.0179047f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_331 N_A_M1031_g N_A_604_419#_c_1123_n 0.00683691f $X=3.915 $Y=2.415 $X2=0
+ $Y2=0
cc_332 N_A_c_205_n N_A_604_419#_c_1123_n 0.0176376f $X=3.99 $Y=1.65 $X2=0 $Y2=0
cc_333 N_A_M1030_g N_A_37_131#_c_1272_n 0.0156733f $X=0.525 $Y=0.865 $X2=0 $Y2=0
cc_334 N_A_c_196_n N_A_37_131#_c_1272_n 0.0228597f $X=0.425 $Y=1.535 $X2=0 $Y2=0
cc_335 N_A_c_197_n N_A_37_131#_c_1272_n 0.00123254f $X=0.425 $Y=1.535 $X2=0
+ $Y2=0
cc_336 N_A_c_196_n N_A_37_131#_c_1273_n 0.0124839f $X=0.425 $Y=1.535 $X2=0 $Y2=0
cc_337 N_A_c_197_n N_A_37_131#_c_1273_n 0.00404657f $X=0.425 $Y=1.535 $X2=0
+ $Y2=0
cc_338 N_A_M1030_g N_A_37_131#_c_1274_n 7.169e-19 $X=0.525 $Y=0.865 $X2=0 $Y2=0
cc_339 N_A_M1030_g N_VGND_c_1297_n 0.0122088f $X=0.525 $Y=0.865 $X2=0 $Y2=0
cc_340 N_A_M1016_g N_VGND_c_1298_n 0.00930558f $X=2.355 $Y=0.865 $X2=0 $Y2=0
cc_341 N_A_c_198_n N_VGND_c_1298_n 0.00373826f $X=2.38 $Y=1.915 $X2=0 $Y2=0
cc_342 N_A_c_202_n N_VGND_c_1298_n 0.00212447f $X=2.445 $Y=1.43 $X2=0 $Y2=0
cc_343 N_A_c_203_n N_VGND_c_1298_n 0.00640889f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_344 N_A_M1035_g N_VGND_c_1299_n 0.00774903f $X=3.915 $Y=0.865 $X2=0 $Y2=0
cc_345 N_A_M1003_g N_VGND_c_1306_n 0.00313222f $X=5.535 $Y=0.865 $X2=0 $Y2=0
cc_346 N_A_M1030_g N_VGND_c_1312_n 0.00332367f $X=0.525 $Y=0.865 $X2=0 $Y2=0
cc_347 N_A_M1030_g N_VGND_c_1321_n 0.00387424f $X=0.525 $Y=0.865 $X2=0 $Y2=0
cc_348 N_A_M1016_g N_VGND_c_1321_n 8.90604e-19 $X=2.355 $Y=0.865 $X2=0 $Y2=0
cc_349 N_A_M1035_g N_VGND_c_1321_n 9.15004e-19 $X=3.915 $Y=0.865 $X2=0 $Y2=0
cc_350 N_A_M1003_g N_VGND_c_1321_n 0.0046122f $X=5.535 $Y=0.865 $X2=0 $Y2=0
cc_351 N_A_M1035_g N_A_604_131#_c_1435_n 0.0143894f $X=3.915 $Y=0.865 $X2=0
+ $Y2=0
cc_352 N_A_c_220_n N_A_604_131#_c_1435_n 0.00339889f $X=4.825 $Y=1.83 $X2=0
+ $Y2=0
cc_353 N_A_c_203_n N_A_604_131#_c_1435_n 0.0442922f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_354 N_A_c_204_n N_A_604_131#_c_1435_n 7.77126e-19 $X=3.825 $Y=1.77 $X2=0
+ $Y2=0
cc_355 N_A_c_203_n N_A_604_131#_c_1436_n 0.0144739f $X=3.725 $Y=1.65 $X2=0 $Y2=0
cc_356 N_A_328_131#_c_427_n N_CIN_M1025_g 0.00680672f $X=1.78 $Y=0.93 $X2=0
+ $Y2=0
cc_357 N_A_328_131#_c_420_n N_CIN_M1025_g 0.00246631f $X=1.977 $Y=2.192 $X2=0
+ $Y2=0
cc_358 N_A_328_131#_c_405_n N_CIN_M1025_g 0.00213756f $X=1.977 $Y=2.055 $X2=0
+ $Y2=0
cc_359 N_A_328_131#_c_407_n N_CIN_M1025_g 0.00550234f $X=1.825 $Y=1.295 $X2=0
+ $Y2=0
cc_360 N_A_328_131#_c_410_n N_CIN_M1025_g 0.00586343f $X=1.68 $Y=1.295 $X2=0
+ $Y2=0
cc_361 N_A_328_131#_c_427_n N_CIN_c_598_n 4.86113e-19 $X=1.78 $Y=0.93 $X2=0
+ $Y2=0
cc_362 N_A_328_131#_c_406_n N_CIN_M1032_g 0.0101533f $X=4.415 $Y=1.295 $X2=0
+ $Y2=0
cc_363 N_A_328_131#_M1039_g N_CIN_c_600_n 0.00912852f $X=4.345 $Y=0.865 $X2=0
+ $Y2=0
cc_364 N_A_328_131#_M1039_g N_CIN_M1001_g 0.0169417f $X=4.345 $Y=0.865 $X2=0
+ $Y2=0
cc_365 N_A_328_131#_M1012_g N_CIN_M1001_g 0.0239556f $X=4.345 $Y=2.415 $X2=0
+ $Y2=0
cc_366 N_A_328_131#_c_404_n N_CIN_M1001_g 0.0201591f $X=4.365 $Y=1.48 $X2=0
+ $Y2=0
cc_367 N_A_328_131#_c_408_n N_CIN_M1001_g 0.00394929f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_368 N_A_328_131#_c_409_n N_CIN_M1001_g 0.00150133f $X=4.705 $Y=1.295 $X2=0
+ $Y2=0
cc_369 N_A_328_131#_c_411_n N_CIN_M1001_g 0.00411222f $X=4.56 $Y=1.295 $X2=0
+ $Y2=0
cc_370 N_A_328_131#_c_427_n CIN 0.0231376f $X=1.78 $Y=0.93 $X2=0 $Y2=0
cc_371 N_A_328_131#_c_406_n CIN 0.00586195f $X=4.415 $Y=1.295 $X2=0 $Y2=0
cc_372 N_A_328_131#_c_407_n CIN 0.00263375f $X=1.825 $Y=1.295 $X2=0 $Y2=0
cc_373 N_A_328_131#_c_410_n CIN 0.0043436f $X=1.68 $Y=1.295 $X2=0 $Y2=0
cc_374 N_A_328_131#_c_407_n N_B_M1005_g 8.80992e-19 $X=1.825 $Y=1.295 $X2=0
+ $Y2=0
cc_375 N_A_328_131#_c_410_n N_B_M1005_g 0.00117948f $X=1.68 $Y=1.295 $X2=0 $Y2=0
cc_376 N_A_328_131#_c_427_n N_B_M1028_g 0.00855994f $X=1.78 $Y=0.93 $X2=0 $Y2=0
cc_377 N_A_328_131#_c_405_n N_B_M1028_g 0.011011f $X=1.977 $Y=2.055 $X2=0 $Y2=0
cc_378 N_A_328_131#_c_407_n N_B_M1028_g 4.82614e-19 $X=1.825 $Y=1.295 $X2=0
+ $Y2=0
cc_379 N_A_328_131#_c_410_n N_B_M1028_g 0.00901048f $X=1.68 $Y=1.295 $X2=0 $Y2=0
cc_380 N_A_328_131#_c_420_n N_B_M1019_g 0.00177618f $X=1.977 $Y=2.192 $X2=0
+ $Y2=0
cc_381 N_A_328_131#_c_429_n N_B_M1019_g 0.00651442f $X=1.935 $Y=2.22 $X2=0 $Y2=0
cc_382 N_A_328_131#_c_405_n N_B_M1019_g 7.69674e-19 $X=1.977 $Y=2.055 $X2=0
+ $Y2=0
cc_383 N_A_328_131#_c_406_n N_B_M1033_g 0.00536679f $X=4.415 $Y=1.295 $X2=0
+ $Y2=0
cc_384 N_A_328_131#_M1012_g N_B_c_702_n 0.0104164f $X=4.345 $Y=2.415 $X2=0 $Y2=0
cc_385 N_A_328_131#_c_408_n N_B_M1008_g 0.00270976f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_386 N_A_328_131#_c_420_n N_B_c_704_n 0.00189002f $X=1.977 $Y=2.192 $X2=0
+ $Y2=0
cc_387 N_A_328_131#_c_405_n N_B_c_704_n 0.00950644f $X=1.977 $Y=2.055 $X2=0
+ $Y2=0
cc_388 N_A_328_131#_c_406_n N_B_c_704_n 0.00259304f $X=4.415 $Y=1.295 $X2=0
+ $Y2=0
cc_389 N_A_328_131#_c_410_n N_B_c_704_n 5.49155e-19 $X=1.68 $Y=1.295 $X2=0 $Y2=0
cc_390 N_A_328_131#_c_405_n B 0.0163782f $X=1.977 $Y=2.055 $X2=0 $Y2=0
cc_391 N_A_328_131#_c_407_n B 0.00750019f $X=1.825 $Y=1.295 $X2=0 $Y2=0
cc_392 N_A_328_131#_c_410_n B 0.0118758f $X=1.68 $Y=1.295 $X2=0 $Y2=0
cc_393 N_A_328_131#_c_408_n N_A_884_131#_M1004_g 0.00582539f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_394 N_A_328_131#_c_408_n N_A_884_131#_M1017_g 0.00290083f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_395 N_A_328_131#_c_408_n N_A_884_131#_M1018_g 0.00290083f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_396 N_A_328_131#_c_395_n N_A_884_131#_M1021_g 0.0160013f $X=7.83 $Y=1.185
+ $X2=0 $Y2=0
cc_397 N_A_328_131#_c_413_n N_A_884_131#_M1021_g 4.30063e-19 $X=8.93 $Y=1.35
+ $X2=0 $Y2=0
cc_398 N_A_328_131#_c_414_n N_A_884_131#_M1021_g 0.0157377f $X=9.12 $Y=1.35
+ $X2=0 $Y2=0
cc_399 N_A_328_131#_c_408_n N_A_884_131#_c_842_n 0.0358306f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_400 N_A_328_131#_c_409_n N_A_884_131#_c_842_n 0.00718101f $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_401 N_A_328_131#_c_411_n N_A_884_131#_c_842_n 0.0109429f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_402 N_A_328_131#_c_408_n N_A_884_131#_c_830_n 0.0278938f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_403 N_A_328_131#_c_408_n N_A_884_131#_c_872_n 0.0282217f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_404 N_A_328_131#_M1012_g N_A_884_131#_c_839_n 2.58065e-19 $X=4.345 $Y=2.415
+ $X2=0 $Y2=0
cc_405 N_A_328_131#_M1010_g N_A_884_131#_c_833_n 0.0256762f $X=7.83 $Y=2.465
+ $X2=0 $Y2=0
cc_406 N_A_328_131#_c_408_n N_A_884_131#_c_833_n 0.0144682f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_407 N_A_328_131#_M1010_g N_VPWR_c_986_n 0.0144704f $X=7.83 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_A_328_131#_M1022_g N_VPWR_c_986_n 7.24342e-19 $X=8.26 $Y=2.465 $X2=0
+ $Y2=0
cc_409 N_A_328_131#_c_413_n N_VPWR_c_986_n 8.03939e-19 $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_410 N_A_328_131#_M1010_g N_VPWR_c_987_n 7.24342e-19 $X=7.83 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A_328_131#_M1022_g N_VPWR_c_987_n 0.0141881f $X=8.26 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A_328_131#_M1023_g N_VPWR_c_987_n 0.0141881f $X=8.69 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A_328_131#_M1037_g N_VPWR_c_987_n 7.24342e-19 $X=9.12 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_A_328_131#_M1023_g N_VPWR_c_989_n 7.24342e-19 $X=8.69 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_A_328_131#_M1037_g N_VPWR_c_989_n 0.0152928f $X=9.12 $Y=2.465 $X2=0
+ $Y2=0
cc_416 N_A_328_131#_M1010_g N_VPWR_c_999_n 0.00486043f $X=7.83 $Y=2.465 $X2=0
+ $Y2=0
cc_417 N_A_328_131#_M1022_g N_VPWR_c_999_n 0.00486043f $X=8.26 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A_328_131#_M1023_g N_VPWR_c_1000_n 0.00486043f $X=8.69 $Y=2.465 $X2=0
+ $Y2=0
cc_419 N_A_328_131#_M1037_g N_VPWR_c_1000_n 0.00486043f $X=9.12 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_A_328_131#_M1012_g N_VPWR_c_980_n 9.39239e-19 $X=4.345 $Y=2.415 $X2=0
+ $Y2=0
cc_421 N_A_328_131#_M1010_g N_VPWR_c_980_n 0.00824727f $X=7.83 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_328_131#_M1022_g N_VPWR_c_980_n 0.00824727f $X=8.26 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_328_131#_M1023_g N_VPWR_c_980_n 0.00824727f $X=8.69 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_328_131#_M1037_g N_VPWR_c_980_n 0.00824727f $X=9.12 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_328_131#_M1012_g N_A_604_419#_c_1123_n 2.38308e-19 $X=4.345 $Y=2.415
+ $X2=0 $Y2=0
cc_426 N_A_328_131#_c_408_n N_SUM_c_1149_n 0.0195745f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_427 N_A_328_131#_c_408_n N_SUM_c_1150_n 0.00608116f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_428 N_A_328_131#_c_408_n N_SUM_c_1153_n 0.0020921f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_429 N_A_328_131#_c_395_n N_SUM_c_1151_n 0.00370118f $X=7.83 $Y=1.185 $X2=0
+ $Y2=0
cc_430 N_A_328_131#_c_408_n N_SUM_c_1151_n 0.0212742f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_431 N_A_328_131#_c_412_n N_SUM_c_1151_n 3.4335e-19 $X=7.92 $Y=1.295 $X2=0
+ $Y2=0
cc_432 N_A_328_131#_c_413_n N_SUM_c_1151_n 0.0035813f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_433 N_A_328_131#_M1010_g SUM 0.00748769f $X=7.83 $Y=2.465 $X2=0 $Y2=0
cc_434 N_A_328_131#_c_408_n SUM 0.0316544f $X=7.775 $Y=1.295 $X2=0 $Y2=0
cc_435 N_A_328_131#_c_412_n SUM 3.32075e-19 $X=7.92 $Y=1.295 $X2=0 $Y2=0
cc_436 N_A_328_131#_c_413_n SUM 0.0219618f $X=8.93 $Y=1.35 $X2=0 $Y2=0
cc_437 N_A_328_131#_c_414_n SUM 9.20478e-19 $X=9.12 $Y=1.35 $X2=0 $Y2=0
cc_438 N_A_328_131#_c_397_n N_COUT_c_1220_n 0.00973732f $X=8.26 $Y=1.185 $X2=0
+ $Y2=0
cc_439 N_A_328_131#_c_399_n N_COUT_c_1220_n 0.00969075f $X=8.69 $Y=1.185 $X2=0
+ $Y2=0
cc_440 N_A_328_131#_c_413_n N_COUT_c_1220_n 0.0428504f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_441 N_A_328_131#_c_414_n N_COUT_c_1220_n 6.95778e-19 $X=9.12 $Y=1.35 $X2=0
+ $Y2=0
cc_442 N_A_328_131#_c_412_n N_COUT_c_1224_n 0.00326755f $X=7.92 $Y=1.295 $X2=0
+ $Y2=0
cc_443 N_A_328_131#_c_413_n N_COUT_c_1224_n 0.0138932f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_444 N_A_328_131#_c_414_n N_COUT_c_1224_n 7.81868e-19 $X=9.12 $Y=1.35 $X2=0
+ $Y2=0
cc_445 N_A_328_131#_M1022_g N_COUT_c_1215_n 0.0134266f $X=8.26 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_A_328_131#_M1023_g N_COUT_c_1215_n 0.0135888f $X=8.69 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_328_131#_c_413_n N_COUT_c_1215_n 0.0377393f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_448 N_A_328_131#_c_414_n N_COUT_c_1215_n 0.00213862f $X=9.12 $Y=1.35 $X2=0
+ $Y2=0
cc_449 N_A_328_131#_M1010_g N_COUT_c_1216_n 9.70174e-19 $X=7.83 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_328_131#_c_412_n N_COUT_c_1216_n 7.75846e-19 $X=7.92 $Y=1.295 $X2=0
+ $Y2=0
cc_451 N_A_328_131#_c_413_n N_COUT_c_1216_n 0.0114721f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_452 N_A_328_131#_c_414_n N_COUT_c_1216_n 0.00224327f $X=9.12 $Y=1.35 $X2=0
+ $Y2=0
cc_453 N_A_328_131#_c_401_n N_COUT_c_1235_n 0.0142044f $X=9.12 $Y=1.185 $X2=0
+ $Y2=0
cc_454 N_A_328_131#_c_413_n N_COUT_c_1235_n 0.0054189f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_455 N_A_328_131#_M1037_g N_COUT_c_1217_n 0.0178269f $X=9.12 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A_328_131#_c_413_n N_COUT_c_1217_n 0.00530126f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_457 N_A_328_131#_c_413_n N_COUT_c_1239_n 0.015412f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_458 N_A_328_131#_c_414_n N_COUT_c_1239_n 7.81868e-19 $X=9.12 $Y=1.35 $X2=0
+ $Y2=0
cc_459 N_A_328_131#_c_413_n N_COUT_c_1218_n 0.0124005f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_460 N_A_328_131#_c_414_n N_COUT_c_1218_n 0.00224327f $X=9.12 $Y=1.35 $X2=0
+ $Y2=0
cc_461 N_A_328_131#_c_401_n COUT 0.0262682f $X=9.12 $Y=1.185 $X2=0 $Y2=0
cc_462 N_A_328_131#_c_413_n COUT 0.0272848f $X=8.93 $Y=1.35 $X2=0 $Y2=0
cc_463 N_A_328_131#_c_427_n N_A_37_131#_c_1274_n 0.0311219f $X=1.78 $Y=0.93
+ $X2=0 $Y2=0
cc_464 N_A_328_131#_c_407_n N_A_37_131#_c_1274_n 0.00153219f $X=1.825 $Y=1.295
+ $X2=0 $Y2=0
cc_465 N_A_328_131#_c_427_n N_VGND_c_1298_n 0.00745143f $X=1.78 $Y=0.93 $X2=0
+ $Y2=0
cc_466 N_A_328_131#_c_406_n N_VGND_c_1298_n 0.00926257f $X=4.415 $Y=1.295 $X2=0
+ $Y2=0
cc_467 N_A_328_131#_c_395_n N_VGND_c_1302_n 0.0110428f $X=7.83 $Y=1.185 $X2=0
+ $Y2=0
cc_468 N_A_328_131#_c_397_n N_VGND_c_1302_n 6.15704e-19 $X=8.26 $Y=1.185 $X2=0
+ $Y2=0
cc_469 N_A_328_131#_c_408_n N_VGND_c_1302_n 0.00840185f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_470 N_A_328_131#_c_413_n N_VGND_c_1302_n 0.00127315f $X=8.93 $Y=1.35 $X2=0
+ $Y2=0
cc_471 N_A_328_131#_c_395_n N_VGND_c_1303_n 5.67328e-19 $X=7.83 $Y=1.185 $X2=0
+ $Y2=0
cc_472 N_A_328_131#_c_397_n N_VGND_c_1303_n 0.00972547f $X=8.26 $Y=1.185 $X2=0
+ $Y2=0
cc_473 N_A_328_131#_c_399_n N_VGND_c_1303_n 0.00972547f $X=8.69 $Y=1.185 $X2=0
+ $Y2=0
cc_474 N_A_328_131#_c_401_n N_VGND_c_1303_n 5.67328e-19 $X=9.12 $Y=1.185 $X2=0
+ $Y2=0
cc_475 N_A_328_131#_c_399_n N_VGND_c_1305_n 5.67328e-19 $X=8.69 $Y=1.185 $X2=0
+ $Y2=0
cc_476 N_A_328_131#_c_401_n N_VGND_c_1305_n 0.0116216f $X=9.12 $Y=1.185 $X2=0
+ $Y2=0
cc_477 N_A_328_131#_c_395_n N_VGND_c_1315_n 0.00486043f $X=7.83 $Y=1.185 $X2=0
+ $Y2=0
cc_478 N_A_328_131#_c_397_n N_VGND_c_1315_n 0.00486043f $X=8.26 $Y=1.185 $X2=0
+ $Y2=0
cc_479 N_A_328_131#_c_399_n N_VGND_c_1316_n 0.00486043f $X=8.69 $Y=1.185 $X2=0
+ $Y2=0
cc_480 N_A_328_131#_c_401_n N_VGND_c_1316_n 0.00486043f $X=9.12 $Y=1.185 $X2=0
+ $Y2=0
cc_481 N_A_328_131#_M1039_g N_VGND_c_1321_n 9.15004e-19 $X=4.345 $Y=0.865 $X2=0
+ $Y2=0
cc_482 N_A_328_131#_c_395_n N_VGND_c_1321_n 0.00824727f $X=7.83 $Y=1.185 $X2=0
+ $Y2=0
cc_483 N_A_328_131#_c_397_n N_VGND_c_1321_n 0.00454119f $X=8.26 $Y=1.185 $X2=0
+ $Y2=0
cc_484 N_A_328_131#_c_399_n N_VGND_c_1321_n 0.00454119f $X=8.69 $Y=1.185 $X2=0
+ $Y2=0
cc_485 N_A_328_131#_c_401_n N_VGND_c_1321_n 0.00454119f $X=9.12 $Y=1.185 $X2=0
+ $Y2=0
cc_486 N_A_328_131#_M1039_g N_A_604_131#_c_1435_n 0.00417478f $X=4.345 $Y=0.865
+ $X2=0 $Y2=0
cc_487 N_A_328_131#_c_403_n N_A_604_131#_c_1435_n 0.00213385f $X=4.475 $Y=1.48
+ $X2=0 $Y2=0
cc_488 N_A_328_131#_c_404_n N_A_604_131#_c_1435_n 6.9883e-19 $X=4.365 $Y=1.48
+ $X2=0 $Y2=0
cc_489 N_A_328_131#_c_406_n N_A_604_131#_c_1435_n 0.0299334f $X=4.415 $Y=1.295
+ $X2=0 $Y2=0
cc_490 N_A_328_131#_c_409_n N_A_604_131#_c_1435_n 0.00143382f $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_491 N_A_328_131#_c_411_n N_A_604_131#_c_1435_n 7.63137e-19 $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_492 N_A_328_131#_c_406_n N_A_604_131#_c_1436_n 0.00655395f $X=4.415 $Y=1.295
+ $X2=0 $Y2=0
cc_493 N_CIN_M1025_g N_B_M1011_g 0.0178513f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_494 N_CIN_M1025_g N_B_M1005_g 0.0242256f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_495 CIN N_B_M1005_g 0.00419874f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_496 N_CIN_M1025_g N_B_c_696_n 0.00978218f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_497 N_CIN_M1025_g N_B_M1028_g 0.0433348f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_498 N_CIN_c_598_n N_B_M1028_g 0.00825049f $X=2.87 $Y=0.21 $X2=0 $Y2=0
cc_499 CIN N_B_M1028_g 0.00893411f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_500 N_CIN_M1025_g N_B_M1019_g 0.0112521f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_501 N_CIN_M1032_g N_B_c_700_n 0.0104164f $X=2.945 $Y=0.865 $X2=0 $Y2=0
cc_502 N_CIN_M1032_g N_B_M1033_g 0.0611247f $X=2.945 $Y=0.865 $X2=0 $Y2=0
cc_503 N_CIN_c_600_n N_B_M1033_g 0.00910836f $X=4.74 $Y=0.21 $X2=0 $Y2=0
cc_504 N_CIN_M1001_g N_B_c_702_n 0.0104164f $X=4.815 $Y=0.865 $X2=0 $Y2=0
cc_505 N_CIN_M1001_g N_B_M1008_g 0.149252f $X=4.815 $Y=0.865 $X2=0 $Y2=0
cc_506 N_CIN_M1025_g N_B_c_704_n 0.00791206f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_507 N_CIN_M1025_g B 0.0123581f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_508 N_CIN_M1025_g N_B_c_694_n 0.0157993f $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_509 N_CIN_c_600_n N_A_884_131#_c_842_n 0.00280426f $X=4.74 $Y=0.21 $X2=0
+ $Y2=0
cc_510 N_CIN_M1001_g N_A_884_131#_c_842_n 0.0138439f $X=4.815 $Y=0.865 $X2=0
+ $Y2=0
cc_511 N_CIN_M1001_g N_A_884_131#_c_846_n 0.011911f $X=4.815 $Y=0.865 $X2=0
+ $Y2=0
cc_512 N_CIN_M1001_g N_A_884_131#_c_839_n 0.00816475f $X=4.815 $Y=0.865 $X2=0
+ $Y2=0
cc_513 N_CIN_M1025_g N_A_27_440#_c_966_n 0.00264366f $X=1.565 $Y=0.865 $X2=0
+ $Y2=0
cc_514 N_CIN_M1025_g N_VPWR_c_981_n 7.48776e-19 $X=1.565 $Y=0.865 $X2=0 $Y2=0
cc_515 N_CIN_M1032_g N_VPWR_c_982_n 0.00165827f $X=2.945 $Y=0.865 $X2=0 $Y2=0
cc_516 N_CIN_M1032_g N_VPWR_c_980_n 9.39239e-19 $X=2.945 $Y=0.865 $X2=0 $Y2=0
cc_517 N_CIN_M1001_g N_VPWR_c_980_n 9.39239e-19 $X=4.815 $Y=0.865 $X2=0 $Y2=0
cc_518 N_CIN_M1032_g N_A_604_419#_c_1122_n 2.38292e-19 $X=2.945 $Y=0.865 $X2=0
+ $Y2=0
cc_519 CIN N_A_37_131#_c_1272_n 3.44177e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_520 N_CIN_M1025_g N_A_37_131#_c_1274_n 0.00362493f $X=1.565 $Y=0.865 $X2=0
+ $Y2=0
cc_521 CIN N_A_37_131#_c_1274_n 0.0245041f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_522 N_CIN_c_604_n N_A_37_131#_c_1274_n 3.55221e-19 $X=1.515 $Y=0.21 $X2=0
+ $Y2=0
cc_523 CIN N_VGND_c_1297_n 0.0324763f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_524 N_CIN_c_604_n N_VGND_c_1297_n 0.00381076f $X=1.515 $Y=0.21 $X2=0 $Y2=0
cc_525 N_CIN_c_598_n N_VGND_c_1298_n 0.027048f $X=2.87 $Y=0.21 $X2=0 $Y2=0
cc_526 N_CIN_M1032_g N_VGND_c_1298_n 0.0187168f $X=2.945 $Y=0.865 $X2=0 $Y2=0
cc_527 CIN N_VGND_c_1298_n 0.0310428f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_528 N_CIN_M1032_g N_VGND_c_1299_n 0.00788152f $X=2.945 $Y=0.865 $X2=0 $Y2=0
cc_529 N_CIN_c_600_n N_VGND_c_1299_n 0.0273725f $X=4.74 $Y=0.21 $X2=0 $Y2=0
cc_530 N_CIN_c_600_n N_VGND_c_1306_n 0.0343003f $X=4.74 $Y=0.21 $X2=0 $Y2=0
cc_531 CIN N_VGND_c_1313_n 0.0721327f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_532 N_CIN_c_604_n N_VGND_c_1313_n 0.0243372f $X=1.515 $Y=0.21 $X2=0 $Y2=0
cc_533 N_CIN_c_598_n N_VGND_c_1314_n 0.0241947f $X=2.87 $Y=0.21 $X2=0 $Y2=0
cc_534 N_CIN_c_598_n N_VGND_c_1321_n 0.0265854f $X=2.87 $Y=0.21 $X2=0 $Y2=0
cc_535 N_CIN_c_600_n N_VGND_c_1321_n 0.0555647f $X=4.74 $Y=0.21 $X2=0 $Y2=0
cc_536 N_CIN_c_602_n N_VGND_c_1321_n 0.00930383f $X=2.945 $Y=0.21 $X2=0 $Y2=0
cc_537 CIN N_VGND_c_1321_n 0.0403938f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_538 N_CIN_c_604_n N_VGND_c_1321_n 0.00986799f $X=1.515 $Y=0.21 $X2=0 $Y2=0
cc_539 N_CIN_c_600_n N_A_604_131#_c_1449_n 0.00396765f $X=4.74 $Y=0.21 $X2=0
+ $Y2=0
cc_540 N_CIN_M1032_g N_A_604_131#_c_1436_n 0.00451277f $X=2.945 $Y=0.865 $X2=0
+ $Y2=0
cc_541 N_CIN_c_600_n N_A_604_131#_c_1451_n 0.00514494f $X=4.74 $Y=0.21 $X2=0
+ $Y2=0
cc_542 N_B_M1008_g N_A_884_131#_c_842_n 0.0162169f $X=5.175 $Y=0.865 $X2=0 $Y2=0
cc_543 N_B_M1008_g N_A_884_131#_c_846_n 0.0153909f $X=5.175 $Y=0.865 $X2=0 $Y2=0
cc_544 N_B_c_702_n N_A_884_131#_c_839_n 0.00629506f $X=5.1 $Y=3.15 $X2=0 $Y2=0
cc_545 N_B_M1008_g N_A_884_131#_c_839_n 0.00240721f $X=5.175 $Y=0.865 $X2=0
+ $Y2=0
cc_546 N_B_M1011_g N_A_27_440#_c_963_n 0.0142305f $X=0.905 $Y=2.52 $X2=0 $Y2=0
cc_547 N_B_c_696_n N_A_27_440#_c_963_n 8.54994e-19 $X=2.075 $Y=3.15 $X2=0 $Y2=0
cc_548 N_B_M1011_g N_A_27_440#_c_966_n 0.00436421f $X=0.905 $Y=2.52 $X2=0 $Y2=0
cc_549 N_B_c_696_n N_A_27_440#_c_966_n 0.00357357f $X=2.075 $Y=3.15 $X2=0 $Y2=0
cc_550 N_B_M1011_g N_VPWR_c_981_n 0.0143695f $X=0.905 $Y=2.52 $X2=0 $Y2=0
cc_551 N_B_c_697_n N_VPWR_c_981_n 0.00763335f $X=0.98 $Y=3.15 $X2=0 $Y2=0
cc_552 N_B_M1019_g N_VPWR_c_982_n 8.00091e-19 $X=2.15 $Y=2.415 $X2=0 $Y2=0
cc_553 N_B_c_700_n N_VPWR_c_982_n 0.0191272f $X=3.3 $Y=3.15 $X2=0 $Y2=0
cc_554 N_B_M1033_g N_VPWR_c_982_n 0.00377553f $X=3.375 $Y=0.865 $X2=0 $Y2=0
cc_555 N_B_M1033_g N_VPWR_c_983_n 0.00817367f $X=3.375 $Y=0.865 $X2=0 $Y2=0
cc_556 N_B_c_702_n N_VPWR_c_983_n 0.0237652f $X=5.1 $Y=3.15 $X2=0 $Y2=0
cc_557 N_B_M1008_g N_VPWR_c_984_n 0.00908152f $X=5.175 $Y=0.865 $X2=0 $Y2=0
cc_558 N_B_c_702_n N_VPWR_c_990_n 0.0449431f $X=5.1 $Y=3.15 $X2=0 $Y2=0
cc_559 N_B_c_697_n N_VPWR_c_997_n 0.0480654f $X=0.98 $Y=3.15 $X2=0 $Y2=0
cc_560 N_B_c_700_n N_VPWR_c_998_n 0.0201606f $X=3.3 $Y=3.15 $X2=0 $Y2=0
cc_561 N_B_c_696_n N_VPWR_c_980_n 0.0366384f $X=2.075 $Y=3.15 $X2=0 $Y2=0
cc_562 N_B_c_697_n N_VPWR_c_980_n 0.00749832f $X=0.98 $Y=3.15 $X2=0 $Y2=0
cc_563 N_B_c_700_n N_VPWR_c_980_n 0.0259979f $X=3.3 $Y=3.15 $X2=0 $Y2=0
cc_564 N_B_c_702_n N_VPWR_c_980_n 0.0575032f $X=5.1 $Y=3.15 $X2=0 $Y2=0
cc_565 N_B_c_705_n N_VPWR_c_980_n 0.00370846f $X=2.15 $Y=3.15 $X2=0 $Y2=0
cc_566 N_B_c_706_n N_VPWR_c_980_n 0.00907872f $X=3.375 $Y=3.15 $X2=0 $Y2=0
cc_567 N_B_M1033_g N_A_604_419#_c_1124_n 0.0133411f $X=3.375 $Y=0.865 $X2=0
+ $Y2=0
cc_568 N_B_c_700_n N_A_604_419#_c_1122_n 0.00374851f $X=3.3 $Y=3.15 $X2=0 $Y2=0
cc_569 N_B_M1033_g N_A_604_419#_c_1122_n 2.45679e-19 $X=3.375 $Y=0.865 $X2=0
+ $Y2=0
cc_570 N_B_M1033_g N_A_604_419#_c_1123_n 6.71015e-19 $X=3.375 $Y=0.865 $X2=0
+ $Y2=0
cc_571 N_B_c_702_n N_A_604_419#_c_1123_n 0.00550623f $X=5.1 $Y=3.15 $X2=0 $Y2=0
cc_572 N_B_M1005_g N_A_37_131#_c_1272_n 0.0123273f $X=1.035 $Y=0.865 $X2=0 $Y2=0
cc_573 B N_A_37_131#_c_1272_n 0.00914253f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_574 N_B_c_694_n N_A_37_131#_c_1272_n 0.00381382f $X=1.04 $Y=1.665 $X2=0 $Y2=0
cc_575 N_B_M1005_g N_A_37_131#_c_1274_n 0.0080054f $X=1.035 $Y=0.865 $X2=0 $Y2=0
cc_576 B N_A_37_131#_c_1274_n 0.0170066f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_577 N_B_c_694_n N_A_37_131#_c_1274_n 0.00211206f $X=1.04 $Y=1.665 $X2=0 $Y2=0
cc_578 N_B_M1005_g N_VGND_c_1297_n 0.00259378f $X=1.035 $Y=0.865 $X2=0 $Y2=0
cc_579 N_B_M1028_g N_VGND_c_1298_n 0.00151472f $X=1.995 $Y=0.865 $X2=0 $Y2=0
cc_580 N_B_M1033_g N_VGND_c_1299_n 0.00662319f $X=3.375 $Y=0.865 $X2=0 $Y2=0
cc_581 N_B_M1008_g N_VGND_c_1306_n 0.00313222f $X=5.175 $Y=0.865 $X2=0 $Y2=0
cc_582 N_B_M1005_g N_VGND_c_1313_n 0.00318453f $X=1.035 $Y=0.865 $X2=0 $Y2=0
cc_583 N_B_M1005_g N_VGND_c_1321_n 0.00353602f $X=1.035 $Y=0.865 $X2=0 $Y2=0
cc_584 N_B_M1033_g N_VGND_c_1321_n 8.90604e-19 $X=3.375 $Y=0.865 $X2=0 $Y2=0
cc_585 N_B_M1008_g N_VGND_c_1321_n 0.0046122f $X=5.175 $Y=0.865 $X2=0 $Y2=0
cc_586 N_B_M1033_g N_A_604_131#_c_1435_n 0.01417f $X=3.375 $Y=0.865 $X2=0 $Y2=0
cc_587 N_A_884_131#_c_846_n N_VPWR_M1029_d 0.0111917f $X=5.89 $Y=2.18 $X2=0
+ $Y2=0
cc_588 N_A_884_131#_c_831_n N_VPWR_M1029_d 0.00327294f $X=5.975 $Y=2.095 $X2=0
+ $Y2=0
cc_589 N_A_884_131#_M1000_g N_VPWR_c_984_n 0.0121833f $X=6.11 $Y=2.465 $X2=0
+ $Y2=0
cc_590 N_A_884_131#_M1013_g N_VPWR_c_984_n 6.30983e-19 $X=6.54 $Y=2.465 $X2=0
+ $Y2=0
cc_591 N_A_884_131#_c_846_n N_VPWR_c_984_n 0.022778f $X=5.89 $Y=2.18 $X2=0 $Y2=0
cc_592 N_A_884_131#_M1000_g N_VPWR_c_985_n 7.24342e-19 $X=6.11 $Y=2.465 $X2=0
+ $Y2=0
cc_593 N_A_884_131#_M1013_g N_VPWR_c_985_n 0.0141881f $X=6.54 $Y=2.465 $X2=0
+ $Y2=0
cc_594 N_A_884_131#_M1020_g N_VPWR_c_985_n 0.0141881f $X=6.97 $Y=2.465 $X2=0
+ $Y2=0
cc_595 N_A_884_131#_M1027_g N_VPWR_c_985_n 7.24342e-19 $X=7.4 $Y=2.465 $X2=0
+ $Y2=0
cc_596 N_A_884_131#_M1020_g N_VPWR_c_986_n 7.24342e-19 $X=6.97 $Y=2.465 $X2=0
+ $Y2=0
cc_597 N_A_884_131#_M1027_g N_VPWR_c_986_n 0.01415f $X=7.4 $Y=2.465 $X2=0 $Y2=0
cc_598 N_A_884_131#_c_839_n N_VPWR_c_990_n 0.00735486f $X=4.58 $Y=2.26 $X2=0
+ $Y2=0
cc_599 N_A_884_131#_M1000_g N_VPWR_c_992_n 0.00486043f $X=6.11 $Y=2.465 $X2=0
+ $Y2=0
cc_600 N_A_884_131#_M1013_g N_VPWR_c_992_n 0.00486043f $X=6.54 $Y=2.465 $X2=0
+ $Y2=0
cc_601 N_A_884_131#_M1020_g N_VPWR_c_994_n 0.00486043f $X=6.97 $Y=2.465 $X2=0
+ $Y2=0
cc_602 N_A_884_131#_M1027_g N_VPWR_c_994_n 0.00486043f $X=7.4 $Y=2.465 $X2=0
+ $Y2=0
cc_603 N_A_884_131#_M1000_g N_VPWR_c_980_n 0.00824727f $X=6.11 $Y=2.465 $X2=0
+ $Y2=0
cc_604 N_A_884_131#_M1013_g N_VPWR_c_980_n 0.00824727f $X=6.54 $Y=2.465 $X2=0
+ $Y2=0
cc_605 N_A_884_131#_M1020_g N_VPWR_c_980_n 0.00824727f $X=6.97 $Y=2.465 $X2=0
+ $Y2=0
cc_606 N_A_884_131#_M1027_g N_VPWR_c_980_n 0.00824727f $X=7.4 $Y=2.465 $X2=0
+ $Y2=0
cc_607 N_A_884_131#_c_839_n N_VPWR_c_980_n 0.00874363f $X=4.58 $Y=2.26 $X2=0
+ $Y2=0
cc_608 N_A_884_131#_c_839_n N_A_604_419#_c_1123_n 0.00237494f $X=4.58 $Y=2.26
+ $X2=0 $Y2=0
cc_609 N_A_884_131#_c_846_n A_978_419# 0.00496486f $X=5.89 $Y=2.18 $X2=-0.19
+ $Y2=-0.245
cc_610 N_A_884_131#_c_846_n A_1050_419# 0.00524328f $X=5.89 $Y=2.18 $X2=-0.19
+ $Y2=-0.245
cc_611 N_A_884_131#_M1017_g N_SUM_c_1149_n 0.0138493f $X=6.54 $Y=0.655 $X2=0
+ $Y2=0
cc_612 N_A_884_131#_M1018_g N_SUM_c_1149_n 0.014155f $X=6.97 $Y=0.655 $X2=0
+ $Y2=0
cc_613 N_A_884_131#_c_872_n N_SUM_c_1149_n 0.0338835f $X=6.88 $Y=1.48 $X2=0
+ $Y2=0
cc_614 N_A_884_131#_c_833_n N_SUM_c_1149_n 0.00196854f $X=7.4 $Y=1.48 $X2=0
+ $Y2=0
cc_615 N_A_884_131#_M1004_g N_SUM_c_1150_n 0.00123338f $X=6.11 $Y=0.655 $X2=0
+ $Y2=0
cc_616 N_A_884_131#_c_830_n N_SUM_c_1150_n 0.0130755f $X=5.975 $Y=1.395 $X2=0
+ $Y2=0
cc_617 N_A_884_131#_c_872_n N_SUM_c_1150_n 0.0120711f $X=6.88 $Y=1.48 $X2=0
+ $Y2=0
cc_618 N_A_884_131#_c_833_n N_SUM_c_1150_n 0.00196569f $X=7.4 $Y=1.48 $X2=0
+ $Y2=0
cc_619 N_A_884_131#_M1013_g N_SUM_c_1153_n 0.0137757f $X=6.54 $Y=2.465 $X2=0
+ $Y2=0
cc_620 N_A_884_131#_M1020_g N_SUM_c_1153_n 0.0139586f $X=6.97 $Y=2.465 $X2=0
+ $Y2=0
cc_621 N_A_884_131#_c_872_n N_SUM_c_1153_n 0.0414104f $X=6.88 $Y=1.48 $X2=0
+ $Y2=0
cc_622 N_A_884_131#_c_833_n N_SUM_c_1153_n 0.00247143f $X=7.4 $Y=1.48 $X2=0
+ $Y2=0
cc_623 N_A_884_131#_M1000_g N_SUM_c_1154_n 8.20937e-19 $X=6.11 $Y=2.465 $X2=0
+ $Y2=0
cc_624 N_A_884_131#_c_831_n N_SUM_c_1154_n 0.0110851f $X=5.975 $Y=2.095 $X2=0
+ $Y2=0
cc_625 N_A_884_131#_c_872_n N_SUM_c_1154_n 0.0143593f $X=6.88 $Y=1.48 $X2=0
+ $Y2=0
cc_626 N_A_884_131#_c_833_n N_SUM_c_1154_n 0.00256759f $X=7.4 $Y=1.48 $X2=0
+ $Y2=0
cc_627 N_A_884_131#_M1021_g N_SUM_c_1151_n 0.0122443f $X=7.4 $Y=0.655 $X2=0
+ $Y2=0
cc_628 N_A_884_131#_c_833_n N_SUM_c_1151_n 0.00189961f $X=7.4 $Y=1.48 $X2=0
+ $Y2=0
cc_629 N_A_884_131#_M1018_g SUM 7.02698e-19 $X=6.97 $Y=0.655 $X2=0 $Y2=0
cc_630 N_A_884_131#_M1020_g SUM 9.54489e-19 $X=6.97 $Y=2.465 $X2=0 $Y2=0
cc_631 N_A_884_131#_M1021_g SUM 0.00258965f $X=7.4 $Y=0.655 $X2=0 $Y2=0
cc_632 N_A_884_131#_M1027_g SUM 0.014474f $X=7.4 $Y=2.465 $X2=0 $Y2=0
cc_633 N_A_884_131#_c_872_n SUM 0.0134955f $X=6.88 $Y=1.48 $X2=0 $Y2=0
cc_634 N_A_884_131#_c_833_n SUM 0.0224148f $X=7.4 $Y=1.48 $X2=0 $Y2=0
cc_635 N_A_884_131#_c_842_n N_VGND_M1003_d 0.00714584f $X=5.89 $Y=0.865 $X2=0
+ $Y2=0
cc_636 N_A_884_131#_c_830_n N_VGND_M1003_d 5.56021e-19 $X=5.975 $Y=1.395 $X2=0
+ $Y2=0
cc_637 N_A_884_131#_M1004_g N_VGND_c_1300_n 0.00700872f $X=6.11 $Y=0.655 $X2=0
+ $Y2=0
cc_638 N_A_884_131#_M1017_g N_VGND_c_1300_n 5.17829e-19 $X=6.54 $Y=0.655 $X2=0
+ $Y2=0
cc_639 N_A_884_131#_c_842_n N_VGND_c_1300_n 0.0224006f $X=5.89 $Y=0.865 $X2=0
+ $Y2=0
cc_640 N_A_884_131#_M1004_g N_VGND_c_1301_n 6.33489e-19 $X=6.11 $Y=0.655 $X2=0
+ $Y2=0
cc_641 N_A_884_131#_M1017_g N_VGND_c_1301_n 0.011104f $X=6.54 $Y=0.655 $X2=0
+ $Y2=0
cc_642 N_A_884_131#_M1018_g N_VGND_c_1301_n 0.0110576f $X=6.97 $Y=0.655 $X2=0
+ $Y2=0
cc_643 N_A_884_131#_M1021_g N_VGND_c_1301_n 6.25324e-19 $X=7.4 $Y=0.655 $X2=0
+ $Y2=0
cc_644 N_A_884_131#_M1018_g N_VGND_c_1302_n 6.25324e-19 $X=6.97 $Y=0.655 $X2=0
+ $Y2=0
cc_645 N_A_884_131#_M1021_g N_VGND_c_1302_n 0.0110098f $X=7.4 $Y=0.655 $X2=0
+ $Y2=0
cc_646 N_A_884_131#_c_842_n N_VGND_c_1306_n 0.0161765f $X=5.89 $Y=0.865 $X2=0
+ $Y2=0
cc_647 N_A_884_131#_M1004_g N_VGND_c_1308_n 0.00544954f $X=6.11 $Y=0.655 $X2=0
+ $Y2=0
cc_648 N_A_884_131#_M1017_g N_VGND_c_1308_n 0.00486043f $X=6.54 $Y=0.655 $X2=0
+ $Y2=0
cc_649 N_A_884_131#_c_842_n N_VGND_c_1308_n 3.02166e-19 $X=5.89 $Y=0.865 $X2=0
+ $Y2=0
cc_650 N_A_884_131#_M1018_g N_VGND_c_1310_n 0.00486043f $X=6.97 $Y=0.655 $X2=0
+ $Y2=0
cc_651 N_A_884_131#_M1021_g N_VGND_c_1310_n 0.00486043f $X=7.4 $Y=0.655 $X2=0
+ $Y2=0
cc_652 N_A_884_131#_M1004_g N_VGND_c_1321_n 0.008811f $X=6.11 $Y=0.655 $X2=0
+ $Y2=0
cc_653 N_A_884_131#_M1017_g N_VGND_c_1321_n 0.00824727f $X=6.54 $Y=0.655 $X2=0
+ $Y2=0
cc_654 N_A_884_131#_M1018_g N_VGND_c_1321_n 0.00824727f $X=6.97 $Y=0.655 $X2=0
+ $Y2=0
cc_655 N_A_884_131#_M1021_g N_VGND_c_1321_n 0.00824727f $X=7.4 $Y=0.655 $X2=0
+ $Y2=0
cc_656 N_A_884_131#_c_842_n N_VGND_c_1321_n 0.03383f $X=5.89 $Y=0.865 $X2=0
+ $Y2=0
cc_657 N_A_884_131#_c_842_n A_978_131# 0.00306022f $X=5.89 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_658 N_A_884_131#_c_842_n A_1050_131# 0.00307396f $X=5.89 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_659 N_A_27_440#_c_963_n N_VPWR_M1038_d 0.00357407f $X=1.11 $Y=2.365 $X2=-0.19
+ $Y2=1.655
cc_660 N_A_27_440#_c_957_n N_VPWR_c_981_n 0.00858833f $X=0.26 $Y=2.685 $X2=0
+ $Y2=0
cc_661 N_A_27_440#_c_963_n N_VPWR_c_981_n 0.0170777f $X=1.11 $Y=2.365 $X2=0
+ $Y2=0
cc_662 N_A_27_440#_c_957_n N_VPWR_c_996_n 0.00722588f $X=0.26 $Y=2.685 $X2=0
+ $Y2=0
cc_663 N_A_27_440#_c_966_n N_VPWR_c_997_n 0.0031876f $X=1.215 $Y=2.365 $X2=0
+ $Y2=0
cc_664 N_A_27_440#_c_957_n N_VPWR_c_980_n 0.00840852f $X=0.26 $Y=2.685 $X2=0
+ $Y2=0
cc_665 N_A_27_440#_c_966_n N_VPWR_c_980_n 0.0049224f $X=1.215 $Y=2.365 $X2=0
+ $Y2=0
cc_666 N_VPWR_M1009_d N_A_604_419#_c_1124_n 0.00593111f $X=3.45 $Y=2.095 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_983_n N_A_604_419#_c_1124_n 0.022455f $X=3.645 $Y=2.56 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_982_n N_A_604_419#_c_1122_n 0.00229149f $X=2.73 $Y=2.27 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_983_n N_A_604_419#_c_1122_n 0.0020718f $X=3.645 $Y=2.56 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_998_n N_A_604_419#_c_1122_n 0.00583743f $X=3.48 $Y=3.33 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_980_n N_A_604_419#_c_1122_n 0.00693148f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_983_n N_A_604_419#_c_1123_n 0.0132812f $X=3.645 $Y=2.56 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_990_n N_A_604_419#_c_1123_n 0.00651952f $X=5.73 $Y=3.33 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_980_n N_A_604_419#_c_1123_n 0.00775969f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_980_n N_SUM_M1000_s 0.00536646f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_676 N_VPWR_c_980_n N_SUM_M1020_s 0.00536646f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_677 N_VPWR_c_992_n N_SUM_c_1194_n 0.0124525f $X=6.59 $Y=3.33 $X2=0 $Y2=0
cc_678 N_VPWR_c_980_n N_SUM_c_1194_n 0.00730901f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_679 N_VPWR_M1013_d N_SUM_c_1153_n 0.00181369f $X=6.615 $Y=1.835 $X2=0 $Y2=0
cc_680 N_VPWR_c_985_n N_SUM_c_1153_n 0.016476f $X=6.755 $Y=2.19 $X2=0 $Y2=0
cc_681 N_VPWR_c_994_n N_SUM_c_1198_n 0.0124525f $X=7.45 $Y=3.33 $X2=0 $Y2=0
cc_682 N_VPWR_c_980_n N_SUM_c_1198_n 0.00730901f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_683 N_VPWR_M1027_d SUM 0.00157044f $X=7.475 $Y=1.835 $X2=0 $Y2=0
cc_684 N_VPWR_c_986_n SUM 0.00561284f $X=7.615 $Y=2.19 $X2=0 $Y2=0
cc_685 N_VPWR_c_980_n N_COUT_M1010_s 0.00536646f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_686 N_VPWR_c_980_n N_COUT_M1023_s 0.00536646f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_687 N_VPWR_c_999_n N_COUT_c_1247_n 0.0124525f $X=8.31 $Y=3.33 $X2=0 $Y2=0
cc_688 N_VPWR_c_980_n N_COUT_c_1247_n 0.00730901f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_689 N_VPWR_M1022_d N_COUT_c_1215_n 0.00180746f $X=8.335 $Y=1.835 $X2=0 $Y2=0
cc_690 N_VPWR_c_987_n N_COUT_c_1215_n 0.0163515f $X=8.475 $Y=2.19 $X2=0 $Y2=0
cc_691 N_VPWR_c_1000_n N_COUT_c_1251_n 0.0124525f $X=9.17 $Y=3.33 $X2=0 $Y2=0
cc_692 N_VPWR_c_980_n N_COUT_c_1251_n 0.00730901f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_693 N_VPWR_M1037_d N_COUT_c_1217_n 0.0027649f $X=9.195 $Y=1.835 $X2=0 $Y2=0
cc_694 N_VPWR_c_989_n N_COUT_c_1217_n 0.0230335f $X=9.335 $Y=2.19 $X2=0 $Y2=0
cc_695 SUM N_COUT_c_1216_n 0.00652871f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_696 N_SUM_c_1149_n N_VGND_M1017_s 0.00176773f $X=7.09 $Y=1.135 $X2=0 $Y2=0
cc_697 N_SUM_c_1151_n N_VGND_M1021_s 8.89729e-19 $X=7.332 $Y=1.135 $X2=0 $Y2=0
cc_698 N_SUM_c_1149_n N_VGND_c_1301_n 0.016047f $X=7.09 $Y=1.135 $X2=0 $Y2=0
cc_699 N_SUM_c_1151_n N_VGND_c_1302_n 0.00553539f $X=7.332 $Y=1.135 $X2=0 $Y2=0
cc_700 N_SUM_c_1207_p N_VGND_c_1308_n 0.0124525f $X=6.325 $Y=0.42 $X2=0 $Y2=0
cc_701 N_SUM_c_1208_p N_VGND_c_1310_n 0.0124525f $X=7.185 $Y=0.42 $X2=0 $Y2=0
cc_702 N_SUM_M1004_d N_VGND_c_1321_n 0.00536646f $X=6.185 $Y=0.235 $X2=0 $Y2=0
cc_703 N_SUM_M1018_d N_VGND_c_1321_n 0.00536646f $X=7.045 $Y=0.235 $X2=0 $Y2=0
cc_704 N_SUM_c_1207_p N_VGND_c_1321_n 0.00730901f $X=6.325 $Y=0.42 $X2=0 $Y2=0
cc_705 N_SUM_c_1208_p N_VGND_c_1321_n 0.00730901f $X=7.185 $Y=0.42 $X2=0 $Y2=0
cc_706 N_COUT_c_1220_n N_VGND_M1015_d 0.00328233f $X=8.81 $Y=0.925 $X2=0 $Y2=0
cc_707 N_COUT_c_1235_n N_VGND_M1036_d 5.837e-19 $X=9.265 $Y=0.925 $X2=0 $Y2=0
cc_708 COUT N_VGND_M1036_d 0.00292842f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_709 COUT N_VGND_M1036_d 0.00103907f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_710 N_COUT_c_1220_n N_VGND_c_1303_n 0.0167019f $X=8.81 $Y=0.925 $X2=0 $Y2=0
cc_711 N_COUT_c_1235_n N_VGND_c_1305_n 0.00274594f $X=9.265 $Y=0.925 $X2=0 $Y2=0
cc_712 COUT N_VGND_c_1305_n 0.020724f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_713 N_COUT_c_1263_p N_VGND_c_1315_n 0.0124525f $X=8.045 $Y=0.42 $X2=0 $Y2=0
cc_714 N_COUT_c_1264_p N_VGND_c_1316_n 0.0124525f $X=8.905 $Y=0.42 $X2=0 $Y2=0
cc_715 N_COUT_M1014_s N_VGND_c_1321_n 0.00408483f $X=7.905 $Y=0.235 $X2=0 $Y2=0
cc_716 N_COUT_M1034_s N_VGND_c_1321_n 0.0028032f $X=8.765 $Y=0.235 $X2=0 $Y2=0
cc_717 N_COUT_c_1263_p N_VGND_c_1321_n 0.00730901f $X=8.045 $Y=0.42 $X2=0 $Y2=0
cc_718 N_COUT_c_1220_n N_VGND_c_1321_n 0.0108944f $X=8.81 $Y=0.925 $X2=0 $Y2=0
cc_719 N_COUT_c_1264_p N_VGND_c_1321_n 0.00730901f $X=8.905 $Y=0.42 $X2=0 $Y2=0
cc_720 N_COUT_c_1235_n N_VGND_c_1321_n 0.00522141f $X=9.265 $Y=0.925 $X2=0 $Y2=0
cc_721 COUT N_VGND_c_1321_n 0.00128539f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_722 N_A_37_131#_c_1272_n N_VGND_M1030_d 0.00267852f $X=1.085 $Y=1.15
+ $X2=-0.19 $Y2=-0.245
cc_723 N_A_37_131#_c_1272_n N_VGND_c_1297_n 0.0208822f $X=1.085 $Y=1.15 $X2=0
+ $Y2=0
cc_724 N_A_37_131#_c_1295_p N_VGND_c_1312_n 0.00314927f $X=0.31 $Y=0.87 $X2=0
+ $Y2=0
cc_725 N_A_37_131#_c_1295_p N_VGND_c_1321_n 0.0056372f $X=0.31 $Y=0.87 $X2=0
+ $Y2=0
cc_726 N_VGND_c_1321_n N_A_604_131#_c_1449_n 0.00761637f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_727 N_VGND_M1033_d N_A_604_131#_c_1435_n 0.00329873f $X=3.45 $Y=0.655 $X2=0
+ $Y2=0
cc_728 N_VGND_c_1299_n N_A_604_131#_c_1435_n 0.0195827f $X=3.61 $Y=0.78 $X2=0
+ $Y2=0
cc_729 N_VGND_c_1321_n N_A_604_131#_c_1451_n 0.00761637f $X=9.36 $Y=0 $X2=0
+ $Y2=0
