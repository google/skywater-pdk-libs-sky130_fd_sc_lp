* File: sky130_fd_sc_lp__o21ba_2.pxi.spice
* Created: Wed Sep  2 10:16:50 2020
* 
x_PM_SKY130_FD_SC_LP__O21BA_2%B1_N N_B1_N_M1008_g N_B1_N_M1010_g B1_N B1_N
+ N_B1_N_c_71_n PM_SKY130_FD_SC_LP__O21BA_2%B1_N
x_PM_SKY130_FD_SC_LP__O21BA_2%A_186_21# N_A_186_21#_M1007_s N_A_186_21#_M1000_d
+ N_A_186_21#_c_97_n N_A_186_21#_M1001_g N_A_186_21#_c_104_n N_A_186_21#_M1009_g
+ N_A_186_21#_c_98_n N_A_186_21#_M1005_g N_A_186_21#_c_105_n N_A_186_21#_M1011_g
+ N_A_186_21#_c_113_p N_A_186_21#_c_99_n N_A_186_21#_c_155_p N_A_186_21#_c_100_n
+ N_A_186_21#_c_140_p N_A_186_21#_c_101_n N_A_186_21#_c_102_n
+ N_A_186_21#_c_103_n PM_SKY130_FD_SC_LP__O21BA_2%A_186_21#
x_PM_SKY130_FD_SC_LP__O21BA_2%A_28_131# N_A_28_131#_M1008_s N_A_28_131#_M1010_s
+ N_A_28_131#_M1000_g N_A_28_131#_M1007_g N_A_28_131#_c_180_n
+ N_A_28_131#_c_181_n N_A_28_131#_c_175_n N_A_28_131#_c_182_n
+ N_A_28_131#_c_176_n N_A_28_131#_c_177_n N_A_28_131#_c_178_n
+ PM_SKY130_FD_SC_LP__O21BA_2%A_28_131#
x_PM_SKY130_FD_SC_LP__O21BA_2%A2 N_A2_M1006_g N_A2_M1002_g A2 A2 A2 A2
+ N_A2_c_244_n PM_SKY130_FD_SC_LP__O21BA_2%A2
x_PM_SKY130_FD_SC_LP__O21BA_2%A1 N_A1_M1004_g N_A1_M1003_g A1 A1 N_A1_c_281_n
+ PM_SKY130_FD_SC_LP__O21BA_2%A1
x_PM_SKY130_FD_SC_LP__O21BA_2%VPWR N_VPWR_M1010_d N_VPWR_M1011_d N_VPWR_M1004_d
+ N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n
+ N_VPWR_c_309_n VPWR N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_312_n
+ N_VPWR_c_303_n PM_SKY130_FD_SC_LP__O21BA_2%VPWR
x_PM_SKY130_FD_SC_LP__O21BA_2%X N_X_M1001_d N_X_M1009_s N_X_c_352_n X X X X X
+ N_X_c_347_n N_X_c_345_n PM_SKY130_FD_SC_LP__O21BA_2%X
x_PM_SKY130_FD_SC_LP__O21BA_2%VGND N_VGND_M1008_d N_VGND_M1005_s N_VGND_M1002_d
+ N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n VGND N_VGND_c_381_n
+ N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n
+ N_VGND_c_387_n N_VGND_c_388_n PM_SKY130_FD_SC_LP__O21BA_2%VGND
x_PM_SKY130_FD_SC_LP__O21BA_2%A_492_47# N_A_492_47#_M1007_d N_A_492_47#_M1003_d
+ N_A_492_47#_c_441_n N_A_492_47#_c_444_n N_A_492_47#_c_440_n
+ N_A_492_47#_c_437_n N_A_492_47#_c_438_n PM_SKY130_FD_SC_LP__O21BA_2%A_492_47#
cc_1 VNB N_B1_N_M1008_g 0.023091f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.865
cc_2 VNB N_B1_N_M1010_g 0.00624234f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.045
cc_3 VNB B1_N 0.00685146f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_B1_N_c_71_n 0.0333599f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.375
cc_5 VNB N_A_186_21#_c_97_n 0.0189367f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.045
cc_6 VNB N_A_186_21#_c_98_n 0.0191095f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.375
cc_7 VNB N_A_186_21#_c_99_n 0.0140142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_186_21#_c_100_n 0.00806045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_186_21#_c_101_n 0.00415359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_186_21#_c_102_n 0.0042742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_186_21#_c_103_n 0.0719729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_28_131#_M1007_g 0.0281101f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.375
cc_13 VNB N_A_28_131#_c_175_n 0.0134592f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_14 VNB N_A_28_131#_c_176_n 0.0294706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_28_131#_c_177_n 0.0024194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_28_131#_c_178_n 0.0350491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_M1006_g 0.00608905f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.865
cc_18 VNB N_A2_M1002_g 0.0187528f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.045
cc_19 VNB A2 0.00680749f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A2_c_244_n 0.0341513f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.295
cc_21 VNB N_A1_M1004_g 0.0077487f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.865
cc_22 VNB N_A1_M1003_g 0.0249327f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.045
cc_23 VNB A1 0.0216363f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_24 VNB N_A1_c_281_n 0.0422969f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.375
cc_25 VNB N_VPWR_c_303_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_345_n 6.33125e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_378_n 0.0163977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_379_n 0.00854837f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.295
cc_29 VNB N_VGND_c_380_n 0.00284395f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_30 VNB N_VGND_c_381_n 0.0179412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_382_n 0.0152106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_383_n 0.029104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_384_n 0.0161295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_385_n 0.224765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_386_n 0.00701736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_387_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_388_n 0.00515832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_492_47#_c_437_n 0.0149276f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.375
cc_39 VNB N_A_492_47#_c_438_n 0.01479f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.54
cc_40 VPB N_B1_N_M1010_g 0.0239243f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.045
cc_41 VPB B1_N 0.00535418f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_42 VPB N_A_186_21#_c_104_n 0.0182421f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_43 VPB N_A_186_21#_c_105_n 0.0176466f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.21
cc_44 VPB N_A_186_21#_c_102_n 0.00307987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_186_21#_c_103_n 0.0206913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_28_131#_M1000_g 0.0200309f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_47 VPB N_A_28_131#_c_180_n 0.0158617f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.54
cc_48 VPB N_A_28_131#_c_181_n 0.00163053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_28_131#_c_182_n 0.0480922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_28_131#_c_176_n 0.0133647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_28_131#_c_178_n 0.00792945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A2_M1006_g 0.0210669f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.865
cc_53 VPB A2 0.00228301f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_54 VPB N_A1_M1004_g 0.0270382f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.865
cc_55 VPB A1 0.00880496f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_56 VPB N_VPWR_c_304_n 0.0208906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_305_n 0.00502094f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.21
cc_58 VPB N_VPWR_c_306_n 0.0115754f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.295
cc_59 VPB N_VPWR_c_307_n 0.0482054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_308_n 0.0311013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_309_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_310_n 0.0179828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_311_n 0.0340041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_312_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_303_n 0.0793975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_X_c_345_n 0.00115646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 N_B1_N_M1008_g N_A_186_21#_c_97_n 0.0123319f $X=0.48 $Y=0.865 $X2=0 $Y2=0
cc_68 N_B1_N_M1010_g N_A_186_21#_c_104_n 0.0134654f $X=0.645 $Y=2.045 $X2=0
+ $Y2=0
cc_69 B1_N N_A_186_21#_c_103_n 0.00437145f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_B1_N_c_71_n N_A_186_21#_c_103_n 0.0335665f $X=0.555 $Y=1.375 $X2=0 $Y2=0
cc_71 N_B1_N_M1010_g N_A_28_131#_c_180_n 0.00822136f $X=0.645 $Y=2.045 $X2=0
+ $Y2=0
cc_72 B1_N N_A_28_131#_c_180_n 0.0100648f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_73 N_B1_N_M1010_g N_A_28_131#_c_182_n 0.0113846f $X=0.645 $Y=2.045 $X2=0
+ $Y2=0
cc_74 B1_N N_A_28_131#_c_182_n 0.010895f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_B1_N_c_71_n N_A_28_131#_c_182_n 0.00236452f $X=0.555 $Y=1.375 $X2=0
+ $Y2=0
cc_76 N_B1_N_M1008_g N_A_28_131#_c_176_n 0.00576874f $X=0.48 $Y=0.865 $X2=0
+ $Y2=0
cc_77 N_B1_N_M1010_g N_A_28_131#_c_176_n 0.0057482f $X=0.645 $Y=2.045 $X2=0
+ $Y2=0
cc_78 B1_N N_A_28_131#_c_176_n 0.0427703f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B1_N_c_71_n N_A_28_131#_c_176_n 0.00786357f $X=0.555 $Y=1.375 $X2=0
+ $Y2=0
cc_80 N_B1_N_M1010_g N_X_c_347_n 0.00347251f $X=0.645 $Y=2.045 $X2=0 $Y2=0
cc_81 N_B1_N_M1008_g N_X_c_345_n 8.90334e-19 $X=0.48 $Y=0.865 $X2=0 $Y2=0
cc_82 N_B1_N_M1010_g N_X_c_345_n 0.0020191f $X=0.645 $Y=2.045 $X2=0 $Y2=0
cc_83 B1_N N_X_c_345_n 0.0431018f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B1_N_c_71_n N_X_c_345_n 3.82667e-19 $X=0.555 $Y=1.375 $X2=0 $Y2=0
cc_85 N_B1_N_M1008_g N_VGND_c_378_n 0.0142412f $X=0.48 $Y=0.865 $X2=0 $Y2=0
cc_86 B1_N N_VGND_c_378_n 0.0283371f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_B1_N_c_71_n N_VGND_c_378_n 0.00111902f $X=0.555 $Y=1.375 $X2=0 $Y2=0
cc_88 N_B1_N_M1008_g N_VGND_c_381_n 0.00332367f $X=0.48 $Y=0.865 $X2=0 $Y2=0
cc_89 N_B1_N_M1008_g N_VGND_c_385_n 0.00387424f $X=0.48 $Y=0.865 $X2=0 $Y2=0
cc_90 N_A_186_21#_c_103_n N_A_28_131#_M1000_g 0.0350034f $X=1.72 $Y=1.455 $X2=0
+ $Y2=0
cc_91 N_A_186_21#_c_113_p N_A_28_131#_M1007_g 7.58189e-19 $X=1.63 $Y=1.35 $X2=0
+ $Y2=0
cc_92 N_A_186_21#_c_101_n N_A_28_131#_M1007_g 0.0172454f $X=2.525 $Y=1.09 $X2=0
+ $Y2=0
cc_93 N_A_186_21#_c_102_n N_A_28_131#_M1007_g 0.00457663f $X=2.51 $Y=1.855 $X2=0
+ $Y2=0
cc_94 N_A_186_21#_c_103_n N_A_28_131#_M1007_g 0.00344571f $X=1.72 $Y=1.455 $X2=0
+ $Y2=0
cc_95 N_A_186_21#_c_104_n N_A_28_131#_c_180_n 0.0156885f $X=1.29 $Y=1.725 $X2=0
+ $Y2=0
cc_96 N_A_186_21#_c_105_n N_A_28_131#_c_180_n 0.0196003f $X=1.72 $Y=1.725 $X2=0
+ $Y2=0
cc_97 N_A_186_21#_c_103_n N_A_28_131#_c_180_n 0.00412679f $X=1.72 $Y=1.455 $X2=0
+ $Y2=0
cc_98 N_A_186_21#_c_102_n N_A_28_131#_c_181_n 0.0109619f $X=2.51 $Y=1.855 $X2=0
+ $Y2=0
cc_99 N_A_186_21#_c_103_n N_A_28_131#_c_181_n 0.0101004f $X=1.72 $Y=1.455 $X2=0
+ $Y2=0
cc_100 N_A_186_21#_c_104_n N_A_28_131#_c_182_n 0.00110351f $X=1.29 $Y=1.725
+ $X2=0 $Y2=0
cc_101 N_A_186_21#_c_113_p N_A_28_131#_c_177_n 0.0105289f $X=1.63 $Y=1.35 $X2=0
+ $Y2=0
cc_102 N_A_186_21#_c_101_n N_A_28_131#_c_177_n 0.020491f $X=2.525 $Y=1.09 $X2=0
+ $Y2=0
cc_103 N_A_186_21#_c_102_n N_A_28_131#_c_177_n 0.0238981f $X=2.51 $Y=1.855 $X2=0
+ $Y2=0
cc_104 N_A_186_21#_c_103_n N_A_28_131#_c_177_n 0.00192158f $X=1.72 $Y=1.455
+ $X2=0 $Y2=0
cc_105 N_A_186_21#_c_113_p N_A_28_131#_c_178_n 6.26417e-19 $X=1.63 $Y=1.35 $X2=0
+ $Y2=0
cc_106 N_A_186_21#_c_101_n N_A_28_131#_c_178_n 0.00372485f $X=2.525 $Y=1.09
+ $X2=0 $Y2=0
cc_107 N_A_186_21#_c_102_n N_A_28_131#_c_178_n 0.00648495f $X=2.51 $Y=1.855
+ $X2=0 $Y2=0
cc_108 N_A_186_21#_c_103_n N_A_28_131#_c_178_n 0.0224656f $X=1.72 $Y=1.455 $X2=0
+ $Y2=0
cc_109 N_A_186_21#_c_101_n N_A2_M1002_g 0.00488216f $X=2.525 $Y=1.09 $X2=0 $Y2=0
cc_110 N_A_186_21#_c_102_n N_A2_M1002_g 7.69809e-19 $X=2.51 $Y=1.855 $X2=0 $Y2=0
cc_111 N_A_186_21#_c_102_n A2 0.0781502f $X=2.51 $Y=1.855 $X2=0 $Y2=0
cc_112 N_A_186_21#_c_102_n N_A2_c_244_n 0.00488502f $X=2.51 $Y=1.855 $X2=0 $Y2=0
cc_113 N_A_186_21#_c_104_n N_VPWR_c_304_n 0.0167531f $X=1.29 $Y=1.725 $X2=0
+ $Y2=0
cc_114 N_A_186_21#_c_105_n N_VPWR_c_304_n 0.00186189f $X=1.72 $Y=1.725 $X2=0
+ $Y2=0
cc_115 N_A_186_21#_c_105_n N_VPWR_c_305_n 0.00463723f $X=1.72 $Y=1.725 $X2=0
+ $Y2=0
cc_116 N_A_186_21#_c_104_n N_VPWR_c_310_n 0.00486043f $X=1.29 $Y=1.725 $X2=0
+ $Y2=0
cc_117 N_A_186_21#_c_105_n N_VPWR_c_310_n 0.00585385f $X=1.72 $Y=1.725 $X2=0
+ $Y2=0
cc_118 N_A_186_21#_c_140_p N_VPWR_c_311_n 0.0135104f $X=2.52 $Y=2.02 $X2=0 $Y2=0
cc_119 N_A_186_21#_M1000_d N_VPWR_c_303_n 0.00509901f $X=2.38 $Y=1.835 $X2=0
+ $Y2=0
cc_120 N_A_186_21#_c_104_n N_VPWR_c_303_n 0.00835506f $X=1.29 $Y=1.725 $X2=0
+ $Y2=0
cc_121 N_A_186_21#_c_105_n N_VPWR_c_303_n 0.0112138f $X=1.72 $Y=1.725 $X2=0
+ $Y2=0
cc_122 N_A_186_21#_c_140_p N_VPWR_c_303_n 0.008076f $X=2.52 $Y=2.02 $X2=0 $Y2=0
cc_123 N_A_186_21#_c_104_n N_X_c_352_n 0.00412148f $X=1.29 $Y=1.725 $X2=0 $Y2=0
cc_124 N_A_186_21#_c_105_n N_X_c_352_n 0.00464178f $X=1.72 $Y=1.725 $X2=0 $Y2=0
cc_125 N_A_186_21#_c_113_p N_X_c_352_n 0.00722203f $X=1.63 $Y=1.35 $X2=0 $Y2=0
cc_126 N_A_186_21#_c_103_n N_X_c_352_n 0.00343036f $X=1.72 $Y=1.455 $X2=0 $Y2=0
cc_127 N_A_186_21#_c_104_n N_X_c_347_n 0.00707776f $X=1.29 $Y=1.725 $X2=0 $Y2=0
cc_128 N_A_186_21#_c_97_n N_X_c_345_n 0.0125052f $X=1.005 $Y=1.185 $X2=0 $Y2=0
cc_129 N_A_186_21#_c_104_n N_X_c_345_n 0.00430375f $X=1.29 $Y=1.725 $X2=0 $Y2=0
cc_130 N_A_186_21#_c_98_n N_X_c_345_n 0.00132046f $X=1.435 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A_186_21#_c_105_n N_X_c_345_n 6.62081e-19 $X=1.72 $Y=1.725 $X2=0 $Y2=0
cc_132 N_A_186_21#_c_113_p N_X_c_345_n 0.0248273f $X=1.63 $Y=1.35 $X2=0 $Y2=0
cc_133 N_A_186_21#_c_155_p N_X_c_345_n 0.011127f $X=1.795 $Y=1.09 $X2=0 $Y2=0
cc_134 N_A_186_21#_c_103_n N_X_c_345_n 0.0330416f $X=1.72 $Y=1.455 $X2=0 $Y2=0
cc_135 N_A_186_21#_c_155_p N_VGND_M1005_s 0.00228167f $X=1.795 $Y=1.09 $X2=0
+ $Y2=0
cc_136 N_A_186_21#_c_97_n N_VGND_c_378_n 0.00590432f $X=1.005 $Y=1.185 $X2=0
+ $Y2=0
cc_137 N_A_186_21#_c_97_n N_VGND_c_379_n 6.92681e-19 $X=1.005 $Y=1.185 $X2=0
+ $Y2=0
cc_138 N_A_186_21#_c_98_n N_VGND_c_379_n 0.0113758f $X=1.435 $Y=1.185 $X2=0
+ $Y2=0
cc_139 N_A_186_21#_c_99_n N_VGND_c_379_n 0.00156694f $X=2.005 $Y=1.09 $X2=0
+ $Y2=0
cc_140 N_A_186_21#_c_155_p N_VGND_c_379_n 0.0221439f $X=1.795 $Y=1.09 $X2=0
+ $Y2=0
cc_141 N_A_186_21#_c_100_n N_VGND_c_379_n 0.0438698f $X=2.17 $Y=0.42 $X2=0 $Y2=0
cc_142 N_A_186_21#_c_103_n N_VGND_c_379_n 0.00133622f $X=1.72 $Y=1.455 $X2=0
+ $Y2=0
cc_143 N_A_186_21#_c_97_n N_VGND_c_382_n 0.00564131f $X=1.005 $Y=1.185 $X2=0
+ $Y2=0
cc_144 N_A_186_21#_c_98_n N_VGND_c_382_n 0.00486043f $X=1.435 $Y=1.185 $X2=0
+ $Y2=0
cc_145 N_A_186_21#_c_100_n N_VGND_c_383_n 0.0178111f $X=2.17 $Y=0.42 $X2=0 $Y2=0
cc_146 N_A_186_21#_M1007_s N_VGND_c_385_n 0.00371702f $X=2.045 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_186_21#_c_97_n N_VGND_c_385_n 0.0114086f $X=1.005 $Y=1.185 $X2=0
+ $Y2=0
cc_148 N_A_186_21#_c_98_n N_VGND_c_385_n 0.00824727f $X=1.435 $Y=1.185 $X2=0
+ $Y2=0
cc_149 N_A_186_21#_c_100_n N_VGND_c_385_n 0.0100304f $X=2.17 $Y=0.42 $X2=0 $Y2=0
cc_150 N_A_186_21#_c_101_n N_A_492_47#_M1007_d 0.00196239f $X=2.525 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_151 N_A_186_21#_c_101_n N_A_492_47#_c_440_n 0.00970967f $X=2.525 $Y=1.09
+ $X2=0 $Y2=0
cc_152 N_A_28_131#_M1000_g N_A2_M1006_g 0.0108801f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_28_131#_M1007_g N_A2_M1002_g 0.0175789f $X=2.385 $Y=0.655 $X2=0 $Y2=0
cc_154 N_A_28_131#_M1007_g A2 2.2289e-19 $X=2.385 $Y=0.655 $X2=0 $Y2=0
cc_155 N_A_28_131#_M1007_g N_A2_c_244_n 0.0176711f $X=2.385 $Y=0.655 $X2=0 $Y2=0
cc_156 N_A_28_131#_c_178_n N_A2_c_244_n 0.0108801f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A_28_131#_c_180_n N_VPWR_M1010_d 0.00576078f $X=2.005 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_158 N_A_28_131#_c_180_n N_VPWR_M1011_d 0.00991233f $X=2.005 $Y=2.375 $X2=0
+ $Y2=0
cc_159 N_A_28_131#_c_181_n N_VPWR_M1011_d 0.00639458f $X=2.12 $Y=2.29 $X2=0
+ $Y2=0
cc_160 N_A_28_131#_c_180_n N_VPWR_c_304_n 0.0220026f $X=2.005 $Y=2.375 $X2=0
+ $Y2=0
cc_161 N_A_28_131#_M1000_g N_VPWR_c_305_n 0.00814323f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_28_131#_c_180_n N_VPWR_c_305_n 0.0271528f $X=2.005 $Y=2.375 $X2=0
+ $Y2=0
cc_163 N_A_28_131#_M1000_g N_VPWR_c_311_n 0.00585385f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_28_131#_M1000_g N_VPWR_c_303_n 0.0111964f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_28_131#_c_180_n N_X_M1009_s 0.00800253f $X=2.005 $Y=2.375 $X2=0 $Y2=0
cc_166 N_A_28_131#_M1000_g N_X_c_352_n 2.18506e-19 $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_28_131#_c_180_n N_X_c_352_n 0.0176511f $X=2.005 $Y=2.375 $X2=0 $Y2=0
cc_168 N_A_28_131#_c_181_n N_X_c_352_n 0.0126217f $X=2.12 $Y=2.29 $X2=0 $Y2=0
cc_169 N_A_28_131#_c_180_n N_X_c_347_n 0.0150969f $X=2.005 $Y=2.375 $X2=0 $Y2=0
cc_170 N_A_28_131#_c_182_n N_X_c_347_n 0.0076648f $X=0.43 $Y=2.085 $X2=0 $Y2=0
cc_171 N_A_28_131#_c_178_n N_X_c_345_n 4.97204e-19 $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A_28_131#_c_176_n N_VGND_c_378_n 5.13382e-19 $X=0.34 $Y=1.92 $X2=0
+ $Y2=0
cc_173 N_A_28_131#_M1007_g N_VGND_c_379_n 0.00320214f $X=2.385 $Y=0.655 $X2=0
+ $Y2=0
cc_174 N_A_28_131#_c_175_n N_VGND_c_381_n 0.00448622f $X=0.265 $Y=0.865 $X2=0
+ $Y2=0
cc_175 N_A_28_131#_M1007_g N_VGND_c_383_n 0.0054895f $X=2.385 $Y=0.655 $X2=0
+ $Y2=0
cc_176 N_A_28_131#_M1007_g N_VGND_c_385_n 0.0112379f $X=2.385 $Y=0.655 $X2=0
+ $Y2=0
cc_177 N_A_28_131#_c_175_n N_VGND_c_385_n 0.00781068f $X=0.265 $Y=0.865 $X2=0
+ $Y2=0
cc_178 N_A_28_131#_M1007_g N_A_492_47#_c_441_n 0.00444742f $X=2.385 $Y=0.655
+ $X2=0 $Y2=0
cc_179 N_A_28_131#_M1007_g N_A_492_47#_c_440_n 0.00225631f $X=2.385 $Y=0.655
+ $X2=0 $Y2=0
cc_180 N_A2_M1006_g N_A1_M1004_g 0.0398505f $X=2.745 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A2_M1002_g N_A1_M1003_g 0.0305383f $X=2.815 $Y=0.655 $X2=0 $Y2=0
cc_182 A2 A1 0.0439654f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A2_c_244_n A1 2.39572e-19 $X=2.87 $Y=1.375 $X2=0 $Y2=0
cc_184 A2 N_A1_c_281_n 0.0121937f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A2_c_244_n N_A1_c_281_n 0.0206067f $X=2.87 $Y=1.375 $X2=0 $Y2=0
cc_186 N_A2_M1006_g N_VPWR_c_307_n 0.00342668f $X=2.745 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A2_M1006_g N_VPWR_c_311_n 0.00551913f $X=2.745 $Y=2.465 $X2=0 $Y2=0
cc_188 A2 N_VPWR_c_311_n 0.00612843f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A2_M1006_g N_VPWR_c_303_n 0.0102094f $X=2.745 $Y=2.465 $X2=0 $Y2=0
cc_190 A2 N_VPWR_c_303_n 0.0119756f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_191 A2 A_564_367# 0.0142716f $X=3.035 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_192 N_A2_M1002_g N_VGND_c_380_n 0.00441214f $X=2.815 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A2_M1002_g N_VGND_c_383_n 0.00417814f $X=2.815 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A2_M1002_g N_VGND_c_385_n 0.00598453f $X=2.815 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A2_M1002_g N_A_492_47#_c_441_n 0.00593619f $X=2.815 $Y=0.655 $X2=0
+ $Y2=0
cc_196 N_A2_M1002_g N_A_492_47#_c_444_n 0.0106027f $X=2.815 $Y=0.655 $X2=0 $Y2=0
cc_197 A2 N_A_492_47#_c_444_n 0.0172948f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A2_c_244_n N_A_492_47#_c_444_n 6.8961e-19 $X=2.87 $Y=1.375 $X2=0 $Y2=0
cc_199 N_A2_M1002_g N_A_492_47#_c_440_n 0.00157927f $X=2.815 $Y=0.655 $X2=0
+ $Y2=0
cc_200 N_A2_c_244_n N_A_492_47#_c_440_n 0.00160319f $X=2.87 $Y=1.375 $X2=0 $Y2=0
cc_201 N_A2_M1002_g N_A_492_47#_c_438_n 0.00105179f $X=2.815 $Y=0.655 $X2=0
+ $Y2=0
cc_202 N_A1_M1004_g N_VPWR_c_307_n 0.0230548f $X=3.32 $Y=2.465 $X2=0 $Y2=0
cc_203 A1 N_VPWR_c_307_n 0.0256672f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_204 N_A1_c_281_n N_VPWR_c_307_n 0.0010583f $X=3.47 $Y=1.375 $X2=0 $Y2=0
cc_205 N_A1_M1004_g N_VPWR_c_311_n 0.00544582f $X=3.32 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A1_M1004_g N_VPWR_c_303_n 0.00964249f $X=3.32 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A1_M1003_g N_VGND_c_380_n 0.00766066f $X=3.325 $Y=0.655 $X2=0 $Y2=0
cc_208 N_A1_M1003_g N_VGND_c_384_n 0.00385517f $X=3.325 $Y=0.655 $X2=0 $Y2=0
cc_209 N_A1_M1003_g N_VGND_c_385_n 0.0054027f $X=3.325 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A1_M1003_g N_A_492_47#_c_441_n 3.20508e-19 $X=3.325 $Y=0.655 $X2=0
+ $Y2=0
cc_211 N_A1_M1003_g N_A_492_47#_c_444_n 0.0135194f $X=3.325 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A1_M1003_g N_A_492_47#_c_438_n 0.00779228f $X=3.325 $Y=0.655 $X2=0
+ $Y2=0
cc_213 A1 N_A_492_47#_c_438_n 0.024971f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_214 N_A1_c_281_n N_A_492_47#_c_438_n 0.00168723f $X=3.47 $Y=1.375 $X2=0 $Y2=0
cc_215 N_VPWR_c_303_n N_X_M1009_s 0.0119922f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_M1010_d N_X_c_347_n 0.00497019f $X=0.72 $Y=1.835 $X2=0 $Y2=0
cc_217 N_VPWR_c_303_n A_564_367# 0.00644681f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_218 N_X_c_345_n N_VGND_c_382_n 0.0150063f $X=1.22 $Y=0.42 $X2=0 $Y2=0
cc_219 N_X_M1001_d N_VGND_c_385_n 0.00380103f $X=1.08 $Y=0.235 $X2=0 $Y2=0
cc_220 N_X_c_345_n N_VGND_c_385_n 0.00950443f $X=1.22 $Y=0.42 $X2=0 $Y2=0
cc_221 N_VGND_c_385_n N_A_492_47#_M1007_d 0.00223559f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_222 N_VGND_c_385_n N_A_492_47#_M1003_d 0.00244241f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_383_n N_A_492_47#_c_441_n 0.0187529f $X=2.935 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_385_n N_A_492_47#_c_441_n 0.0123338f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_M1002_d N_A_492_47#_c_444_n 0.00609649f $X=2.89 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_VGND_c_380_n N_A_492_47#_c_444_n 0.0199082f $X=3.1 $Y=0.38 $X2=0 $Y2=0
cc_227 N_VGND_c_383_n N_A_492_47#_c_444_n 0.00235868f $X=2.935 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_384_n N_A_492_47#_c_444_n 0.0017124f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_385_n N_A_492_47#_c_444_n 0.00816064f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_384_n N_A_492_47#_c_437_n 0.0181384f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_c_385_n N_A_492_47#_c_437_n 0.0104192f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_384_n N_A_492_47#_c_438_n 7.21423e-19 $X=3.6 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_385_n N_A_492_47#_c_438_n 0.00155543f $X=3.6 $Y=0 $X2=0 $Y2=0
