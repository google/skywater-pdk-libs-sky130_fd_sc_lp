* File: sky130_fd_sc_lp__a22o_0.pex.spice
* Created: Wed Sep  2 09:22:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22O_0%A_85_155# 1 2 9 12 15 16 17 18 19 20 22 23 25
+ 26 28 32 36
c87 17 0 1.39434e-19 $X=0.59 $Y=1.445
r88 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=0.94 $X2=0.59 $Y2=0.94
r89 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.925 $Y=2.325
+ $X2=1.925 $Y2=2.63
r90 26 28 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.215 $Y=0.445
+ $X2=1.675 $Y2=0.445
r91 24 26 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.13 $Y=0.61
+ $X2=1.215 $Y2=0.445
r92 24 25 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.13 $Y=0.61
+ $X2=1.13 $Y2=0.775
r93 22 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.76 $Y=2.24
+ $X2=1.925 $Y2=2.325
r94 22 23 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.76 $Y=2.24 $X2=0.76
+ $Y2=2.24
r95 21 35 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.76 $Y=0.86
+ $X2=0.632 $Y2=0.86
r96 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.045 $Y=0.86
+ $X2=1.13 $Y2=0.775
r97 20 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.045 $Y=0.86
+ $X2=0.76 $Y2=0.86
r98 19 23 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.632 $Y=2.155
+ $X2=0.76 $Y2=2.24
r99 18 35 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.632 $Y=0.945
+ $X2=0.632 $Y2=0.86
r100 18 19 54.6846 $w=2.53e-07 $l=1.21e-06 $layer=LI1_cond $X=0.632 $Y=0.945
+ $X2=0.632 $Y2=2.155
r101 16 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=1.28
+ $X2=0.59 $Y2=0.94
r102 16 17 43.0552 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.28
+ $X2=0.59 $Y2=1.445
r103 15 36 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=0.775
+ $X2=0.59 $Y2=0.94
r104 12 17 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=0.66 $Y=2.775
+ $X2=0.66 $Y2=1.445
r105 9 15 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.575 $Y=0.445
+ $X2=0.575 $Y2=0.775
r106 2 32 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=2.455 $X2=1.925 $Y2=2.63
r107 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.675 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%A2 3 7 11 12 13 14 18
c46 13 0 1.39434e-19 $X=1.2 $Y=1.295
r47 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16 $Y=1.5
+ $X2=1.16 $Y2=1.5
r48 14 19 5.20967 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=1.177 $Y=1.665
+ $X2=1.177 $Y2=1.5
r49 13 19 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=1.177 $Y=1.295
+ $X2=1.177 $Y2=1.5
r50 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.84
+ $X2=1.16 $Y2=1.5
r51 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.84
+ $X2=1.16 $Y2=2.005
r52 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.335
+ $X2=1.16 $Y2=1.5
r53 7 12 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.21 $Y=2.775 $X2=1.21
+ $Y2=2.005
r54 3 10 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.1 $Y=0.445 $X2=1.1
+ $Y2=1.335
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%A1 3 6 8 11 13 14 15 16 22 25 29
r46 25 28 88.9594 $w=4.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.9 $Y=1.615
+ $X2=2.9 $Y2=2.12
r47 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.96
+ $Y=1.615 $X2=2.96 $Y2=1.615
r48 15 16 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.035 $Y=1.665
+ $X2=3.035 $Y2=2.035
r49 15 26 1.24592 $w=4.78e-07 $l=5e-08 $layer=LI1_cond $X=3.035 $Y=1.665
+ $X2=3.035 $Y2=1.615
r50 14 26 7.97386 $w=4.78e-07 $l=3.2e-07 $layer=LI1_cond $X=3.035 $Y=1.295
+ $X2=3.035 $Y2=1.615
r51 14 29 6.97712 $w=4.78e-07 $l=2.8e-07 $layer=LI1_cond $X=3.035 $Y=1.295
+ $X2=3.035 $Y2=1.015
r52 13 29 2.60822 $w=4.8e-07 $l=1.18e-07 $layer=LI1_cond $X=3.035 $Y=0.897
+ $X2=3.035 $Y2=1.015
r53 11 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=0.93
+ $X2=1.55 $Y2=0.765
r54 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=0.93 $X2=1.55 $Y2=0.93
r55 8 13 5.30486 $w=2.35e-07 $l=2.4e-07 $layer=LI1_cond $X=2.795 $Y=0.897
+ $X2=3.035 $Y2=0.897
r56 8 10 61.055 $w=2.33e-07 $l=1.245e-06 $layer=LI1_cond $X=2.795 $Y=0.897
+ $X2=1.55 $Y2=0.897
r57 6 28 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.75 $Y=2.775
+ $X2=2.75 $Y2=2.12
r58 3 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.46 $Y=0.445
+ $X2=1.46 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%B1 3 7 12 15 16 17 21
r47 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73 $Y=1.5
+ $X2=1.73 $Y2=1.5
r48 17 22 5.20967 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=1.712 $Y=1.665
+ $X2=1.712 $Y2=1.5
r49 16 22 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=1.712 $Y=1.295
+ $X2=1.712 $Y2=1.5
r50 14 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.73 $Y=1.84
+ $X2=1.73 $Y2=1.5
r51 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.84
+ $X2=1.73 $Y2=2.005
r52 10 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.73 $Y=1.485
+ $X2=1.73 $Y2=1.5
r53 10 12 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.73 $Y=1.41 $X2=2
+ $Y2=1.41
r54 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2 $Y=1.335 $X2=2
+ $Y2=1.41
r55 5 7 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2 $Y=1.335 $X2=2
+ $Y2=0.445
r56 3 15 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.64 $Y=2.775 $X2=1.64
+ $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%B2 3 7 9 10 14
r40 14 17 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.89
+ $X2=2.285 $Y2=2.055
r41 14 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.89
+ $X2=2.285 $Y2=1.725
r42 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=1.89 $X2=2.3 $Y2=1.89
r43 10 15 6.48249 $w=3.98e-07 $l=2.25e-07 $layer=LI1_cond $X=2.265 $Y=1.665
+ $X2=2.265 $Y2=1.89
r44 9 10 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.265 $Y=1.295
+ $X2=2.265 $Y2=1.665
r45 7 16 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=2.36 $Y=0.445
+ $X2=2.36 $Y2=1.725
r46 3 17 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.18 $Y=2.775
+ $X2=2.18 $Y2=2.055
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%X 1 2 7 8 9 10 11 12 13 40 43
r19 43 44 5.7745 $w=5.03e-07 $l=1.15e-07 $layer=LI1_cond $X=0.337 $Y=2.61
+ $X2=0.337 $Y2=2.495
r20 22 35 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=0.595
+ $X2=0.21 $Y2=0.43
r21 13 43 3.90798 $w=5.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.337 $Y=2.775
+ $X2=0.337 $Y2=2.61
r22 12 44 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.21 $Y=2.405 $X2=0.21
+ $Y2=2.495
r23 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=2.035
+ $X2=0.21 $Y2=2.405
r24 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r25 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r26 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=0.925 $X2=0.21
+ $Y2=1.295
r27 7 40 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.24 $Y=0.43 $X2=0.36
+ $Y2=0.43
r28 7 35 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.43 $X2=0.21
+ $Y2=0.43
r29 7 8 14.1981 $w=2.48e-07 $l=3.08e-07 $layer=LI1_cond $X=0.21 $Y=0.617
+ $X2=0.21 $Y2=0.925
r30 7 22 1.01415 $w=2.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.21 $Y=0.617
+ $X2=0.21 $Y2=0.595
r31 2 43 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=2.455 $X2=0.425 $Y2=2.61
r32 1 40 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.235 $X2=0.36 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%VPWR 1 2 9 11 13 16 17 18 24 33
r36 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 24 32 4.36549 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.82 $Y=3.33 $X2=3.09
+ $Y2=3.33
r42 24 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 18 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 16 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=3.33 $X2=0.72
+ $Y2=3.33
r48 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=3.33
+ $X2=0.925 $Y2=3.33
r49 15 26 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.925 $Y2=3.33
r51 11 32 3.2337 $w=3.1e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.975 $Y=3.245
+ $X2=3.09 $Y2=3.33
r52 11 13 23.6065 $w=3.08e-07 $l=6.35e-07 $layer=LI1_cond $X=2.975 $Y=3.245
+ $X2=2.975 $Y2=2.61
r53 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=3.33
r54 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=2.61
r55 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.825
+ $Y=2.455 $X2=2.965 $Y2=2.61
r56 1 9 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=0.735
+ $Y=2.455 $X2=0.925 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%A_257_491# 1 2 9 11 12 15
r24 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.475 $Y=2.905
+ $X2=2.475 $Y2=2.61
r25 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.31 $Y=2.99
+ $X2=2.475 $Y2=2.905
r26 11 12 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.31 $Y=2.99
+ $X2=1.59 $Y2=2.99
r27 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.425 $Y=2.905
+ $X2=1.59 $Y2=2.99
r28 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.425 $Y=2.905
+ $X2=1.425 $Y2=2.61
r29 2 15 300 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_PDIFF $count=2 $X=2.255
+ $Y=2.455 $X2=2.475 $Y2=2.61
r30 1 9 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.285
+ $Y=2.455 $X2=1.425 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__A22O_0%VGND 1 2 11 15 17 19 29 30 33 36
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r46 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.575
+ $Y2=0
r48 27 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=3.12
+ $Y2=0
r49 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r50 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r51 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 22 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r53 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 20 33 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.76
+ $Y2=0
r55 20 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r56 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.575
+ $Y2=0
r57 19 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.16
+ $Y2=0
r58 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r59 17 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r60 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=0.085
+ $X2=2.575 $Y2=0
r61 13 15 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.575 $Y=0.085
+ $X2=2.575 $Y2=0.445
r62 9 33 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0
r63 9 11 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.38
r64 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.235 $X2=2.575 $Y2=0.445
r65 1 11 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.235 $X2=0.79 $Y2=0.38
.ends

